module rain (
    input CLOCK_25,
    input reset,
    input [9:0] h_counter,
    input [9:0] v_counter,
    input [9:0] x_pos,
    input [9:0] y_pos,
    output active_rain
);

reg [32:0] rain_timer;
localparam MAX_TIMER = 200000;


reg rain_draw[95:0][128:0];

always @(posedge CLOCK_25 or posedge reset) begin
    if(reset) begin
        rain_draw[0][0] = 0;rain_draw[1][0] = 0;rain_draw[2][0] = 0;rain_draw[3][0] = 0;rain_draw[4][0] = 0;rain_draw[5][0] = 0;rain_draw[6][0] = 0;rain_draw[7][0] = 0;rain_draw[8][0] = 0;rain_draw[9][0] = 0;rain_draw[10][0] = 0;rain_draw[11][0] = 0;rain_draw[12][0] = 0;rain_draw[13][0] = 0;rain_draw[14][0] = 0;rain_draw[15][0] = 0;rain_draw[16][0] = 0;rain_draw[17][0] = 0;rain_draw[18][0] = 0;rain_draw[19][0] = 0;rain_draw[20][0] = 0;rain_draw[21][0] = 0;rain_draw[22][0] = 0;rain_draw[23][0] = 0;rain_draw[24][0] = 0;rain_draw[25][0] = 0;rain_draw[26][0] = 0;rain_draw[27][0] = 0;rain_draw[28][0] = 0;rain_draw[29][0] = 0;rain_draw[30][0] = 0;rain_draw[31][0] = 0;rain_draw[32][0] = 0;rain_draw[33][0] = 0;rain_draw[34][0] = 0;rain_draw[35][0] = 0;rain_draw[36][0] = 0;rain_draw[37][0] = 0;rain_draw[38][0] = 0;rain_draw[39][0] = 0;rain_draw[40][0] = 0;rain_draw[41][0] = 0;rain_draw[42][0] = 0;rain_draw[43][0] = 0;rain_draw[44][0] = 0;rain_draw[45][0] = 0;rain_draw[46][0] = 0;rain_draw[47][0] = 0;rain_draw[48][0] = 0;rain_draw[49][0] = 0;rain_draw[50][0] = 0;rain_draw[51][0] = 0;rain_draw[52][0] = 0;rain_draw[53][0] = 0;rain_draw[54][0] = 0;rain_draw[55][0] = 0;rain_draw[56][0] = 0;rain_draw[57][0] = 0;rain_draw[58][0] = 0;rain_draw[59][0] = 0;rain_draw[60][0] = 0;rain_draw[61][0] = 0;rain_draw[62][0] = 0;rain_draw[63][0] = 0;rain_draw[64][0] = 0;rain_draw[65][0] = 0;rain_draw[66][0] = 0;rain_draw[67][0] = 0;rain_draw[68][0] = 0;rain_draw[69][0] = 0;rain_draw[70][0] = 0;rain_draw[71][0] = 0;rain_draw[72][0] = 0;rain_draw[73][0] = 0;rain_draw[74][0] = 0;rain_draw[75][0] = 0;rain_draw[76][0] = 0;rain_draw[77][0] = 0;rain_draw[78][0] = 0;rain_draw[79][0] = 0;rain_draw[80][0] = 0;rain_draw[81][0] = 0;rain_draw[82][0] = 0;rain_draw[83][0] = 0;rain_draw[84][0] = 0;rain_draw[85][0] = 0;rain_draw[86][0] = 0;rain_draw[87][0] = 0;rain_draw[88][0] = 0;rain_draw[89][0] = 0;rain_draw[90][0] = 0;rain_draw[91][0] = 0;rain_draw[92][0] = 0;rain_draw[93][0] = 0;rain_draw[94][0] = 0;rain_draw[95][0] = 0;
        rain_draw[0][1] = 0;rain_draw[1][1] = 0;rain_draw[2][1] = 0;rain_draw[3][1] = 0;rain_draw[4][1] = 0;rain_draw[5][1] = 0;rain_draw[6][1] = 0;rain_draw[7][1] = 0;rain_draw[8][1] = 0;rain_draw[9][1] = 0;rain_draw[10][1] = 0;rain_draw[11][1] = 0;rain_draw[12][1] = 0;rain_draw[13][1] = 0;rain_draw[14][1] = 0;rain_draw[15][1] = 0;rain_draw[16][1] = 0;rain_draw[17][1] = 0;rain_draw[18][1] = 0;rain_draw[19][1] = 0;rain_draw[20][1] = 0;rain_draw[21][1] = 0;rain_draw[22][1] = 0;rain_draw[23][1] = 0;rain_draw[24][1] = 0;rain_draw[25][1] = 0;rain_draw[26][1] = 0;rain_draw[27][1] = 0;rain_draw[28][1] = 0;rain_draw[29][1] = 0;rain_draw[30][1] = 0;rain_draw[31][1] = 0;rain_draw[32][1] = 0;rain_draw[33][1] = 0;rain_draw[34][1] = 0;rain_draw[35][1] = 0;rain_draw[36][1] = 0;rain_draw[37][1] = 0;rain_draw[38][1] = 0;rain_draw[39][1] = 0;rain_draw[40][1] = 0;rain_draw[41][1] = 0;rain_draw[42][1] = 0;rain_draw[43][1] = 0;rain_draw[44][1] = 0;rain_draw[45][1] = 0;rain_draw[46][1] = 0;rain_draw[47][1] = 0;rain_draw[48][1] = 0;rain_draw[49][1] = 0;rain_draw[50][1] = 0;rain_draw[51][1] = 0;rain_draw[52][1] = 0;rain_draw[53][1] = 0;rain_draw[54][1] = 0;rain_draw[55][1] = 0;rain_draw[56][1] = 0;rain_draw[57][1] = 0;rain_draw[58][1] = 0;rain_draw[59][1] = 0;rain_draw[60][1] = 0;rain_draw[61][1] = 0;rain_draw[62][1] = 0;rain_draw[63][1] = 0;rain_draw[64][1] = 0;rain_draw[65][1] = 0;rain_draw[66][1] = 0;rain_draw[67][1] = 0;rain_draw[68][1] = 0;rain_draw[69][1] = 0;rain_draw[70][1] = 0;rain_draw[71][1] = 0;rain_draw[72][1] = 0;rain_draw[73][1] = 0;rain_draw[74][1] = 0;rain_draw[75][1] = 0;rain_draw[76][1] = 0;rain_draw[77][1] = 0;rain_draw[78][1] = 0;rain_draw[79][1] = 0;rain_draw[80][1] = 0;rain_draw[81][1] = 0;rain_draw[82][1] = 0;rain_draw[83][1] = 0;rain_draw[84][1] = 0;rain_draw[85][1] = 0;rain_draw[86][1] = 0;rain_draw[87][1] = 0;rain_draw[88][1] = 0;rain_draw[89][1] = 0;rain_draw[90][1] = 0;rain_draw[91][1] = 0;rain_draw[92][1] = 0;rain_draw[93][1] = 0;rain_draw[94][1] = 0;rain_draw[95][1] = 0;
        rain_draw[0][2] = 0;rain_draw[1][2] = 0;rain_draw[2][2] = 0;rain_draw[3][2] = 0;rain_draw[4][2] = 0;rain_draw[5][2] = 0;rain_draw[6][2] = 0;rain_draw[7][2] = 0;rain_draw[8][2] = 0;rain_draw[9][2] = 0;rain_draw[10][2] = 0;rain_draw[11][2] = 0;rain_draw[12][2] = 0;rain_draw[13][2] = 0;rain_draw[14][2] = 0;rain_draw[15][2] = 0;rain_draw[16][2] = 0;rain_draw[17][2] = 0;rain_draw[18][2] = 0;rain_draw[19][2] = 0;rain_draw[20][2] = 0;rain_draw[21][2] = 0;rain_draw[22][2] = 0;rain_draw[23][2] = 0;rain_draw[24][2] = 0;rain_draw[25][2] = 0;rain_draw[26][2] = 0;rain_draw[27][2] = 0;rain_draw[28][2] = 0;rain_draw[29][2] = 0;rain_draw[30][2] = 0;rain_draw[31][2] = 0;rain_draw[32][2] = 0;rain_draw[33][2] = 0;rain_draw[34][2] = 0;rain_draw[35][2] = 0;rain_draw[36][2] = 0;rain_draw[37][2] = 0;rain_draw[38][2] = 0;rain_draw[39][2] = 0;rain_draw[40][2] = 0;rain_draw[41][2] = 0;rain_draw[42][2] = 0;rain_draw[43][2] = 0;rain_draw[44][2] = 0;rain_draw[45][2] = 0;rain_draw[46][2] = 0;rain_draw[47][2] = 0;rain_draw[48][2] = 0;rain_draw[49][2] = 0;rain_draw[50][2] = 0;rain_draw[51][2] = 0;rain_draw[52][2] = 0;rain_draw[53][2] = 0;rain_draw[54][2] = 0;rain_draw[55][2] = 0;rain_draw[56][2] = 0;rain_draw[57][2] = 0;rain_draw[58][2] = 0;rain_draw[59][2] = 0;rain_draw[60][2] = 0;rain_draw[61][2] = 0;rain_draw[62][2] = 0;rain_draw[63][2] = 0;rain_draw[64][2] = 0;rain_draw[65][2] = 0;rain_draw[66][2] = 0;rain_draw[67][2] = 0;rain_draw[68][2] = 0;rain_draw[69][2] = 0;rain_draw[70][2] = 0;rain_draw[71][2] = 0;rain_draw[72][2] = 0;rain_draw[73][2] = 0;rain_draw[74][2] = 0;rain_draw[75][2] = 0;rain_draw[76][2] = 0;rain_draw[77][2] = 0;rain_draw[78][2] = 0;rain_draw[79][2] = 0;rain_draw[80][2] = 0;rain_draw[81][2] = 0;rain_draw[82][2] = 0;rain_draw[83][2] = 0;rain_draw[84][2] = 0;rain_draw[85][2] = 0;rain_draw[86][2] = 0;rain_draw[87][2] = 0;rain_draw[88][2] = 0;rain_draw[89][2] = 0;rain_draw[90][2] = 0;rain_draw[91][2] = 0;rain_draw[92][2] = 0;rain_draw[93][2] = 0;rain_draw[94][2] = 0;rain_draw[95][2] = 0;
        rain_draw[0][3] = 0;rain_draw[1][3] = 0;rain_draw[2][3] = 0;rain_draw[3][3] = 0;rain_draw[4][3] = 0;rain_draw[5][3] = 0;rain_draw[6][3] = 0;rain_draw[7][3] = 0;rain_draw[8][3] = 0;rain_draw[9][3] = 0;rain_draw[10][3] = 0;rain_draw[11][3] = 0;rain_draw[12][3] = 0;rain_draw[13][3] = 0;rain_draw[14][3] = 0;rain_draw[15][3] = 0;rain_draw[16][3] = 0;rain_draw[17][3] = 0;rain_draw[18][3] = 0;rain_draw[19][3] = 0;rain_draw[20][3] = 0;rain_draw[21][3] = 0;rain_draw[22][3] = 0;rain_draw[23][3] = 0;rain_draw[24][3] = 0;rain_draw[25][3] = 0;rain_draw[26][3] = 0;rain_draw[27][3] = 0;rain_draw[28][3] = 0;rain_draw[29][3] = 0;rain_draw[30][3] = 0;rain_draw[31][3] = 0;rain_draw[32][3] = 0;rain_draw[33][3] = 0;rain_draw[34][3] = 0;rain_draw[35][3] = 0;rain_draw[36][3] = 0;rain_draw[37][3] = 0;rain_draw[38][3] = 0;rain_draw[39][3] = 0;rain_draw[40][3] = 0;rain_draw[41][3] = 0;rain_draw[42][3] = 0;rain_draw[43][3] = 0;rain_draw[44][3] = 0;rain_draw[45][3] = 0;rain_draw[46][3] = 0;rain_draw[47][3] = 0;rain_draw[48][3] = 0;rain_draw[49][3] = 0;rain_draw[50][3] = 0;rain_draw[51][3] = 0;rain_draw[52][3] = 0;rain_draw[53][3] = 0;rain_draw[54][3] = 0;rain_draw[55][3] = 0;rain_draw[56][3] = 0;rain_draw[57][3] = 0;rain_draw[58][3] = 0;rain_draw[59][3] = 0;rain_draw[60][3] = 0;rain_draw[61][3] = 0;rain_draw[62][3] = 0;rain_draw[63][3] = 0;rain_draw[64][3] = 0;rain_draw[65][3] = 0;rain_draw[66][3] = 0;rain_draw[67][3] = 0;rain_draw[68][3] = 0;rain_draw[69][3] = 0;rain_draw[70][3] = 0;rain_draw[71][3] = 0;rain_draw[72][3] = 0;rain_draw[73][3] = 0;rain_draw[74][3] = 0;rain_draw[75][3] = 0;rain_draw[76][3] = 0;rain_draw[77][3] = 0;rain_draw[78][3] = 0;rain_draw[79][3] = 0;rain_draw[80][3] = 0;rain_draw[81][3] = 0;rain_draw[82][3] = 0;rain_draw[83][3] = 0;rain_draw[84][3] = 0;rain_draw[85][3] = 0;rain_draw[86][3] = 0;rain_draw[87][3] = 0;rain_draw[88][3] = 0;rain_draw[89][3] = 0;rain_draw[90][3] = 0;rain_draw[91][3] = 0;rain_draw[92][3] = 0;rain_draw[93][3] = 0;rain_draw[94][3] = 0;rain_draw[95][3] = 0;
        rain_draw[0][4] = 0;rain_draw[1][4] = 0;rain_draw[2][4] = 0;rain_draw[3][4] = 0;rain_draw[4][4] = 0;rain_draw[5][4] = 0;rain_draw[6][4] = 0;rain_draw[7][4] = 0;rain_draw[8][4] = 0;rain_draw[9][4] = 0;rain_draw[10][4] = 0;rain_draw[11][4] = 0;rain_draw[12][4] = 0;rain_draw[13][4] = 0;rain_draw[14][4] = 0;rain_draw[15][4] = 0;rain_draw[16][4] = 0;rain_draw[17][4] = 0;rain_draw[18][4] = 0;rain_draw[19][4] = 0;rain_draw[20][4] = 0;rain_draw[21][4] = 0;rain_draw[22][4] = 0;rain_draw[23][4] = 0;rain_draw[24][4] = 0;rain_draw[25][4] = 0;rain_draw[26][4] = 0;rain_draw[27][4] = 0;rain_draw[28][4] = 0;rain_draw[29][4] = 0;rain_draw[30][4] = 0;rain_draw[31][4] = 0;rain_draw[32][4] = 0;rain_draw[33][4] = 0;rain_draw[34][4] = 0;rain_draw[35][4] = 0;rain_draw[36][4] = 0;rain_draw[37][4] = 0;rain_draw[38][4] = 0;rain_draw[39][4] = 0;rain_draw[40][4] = 0;rain_draw[41][4] = 0;rain_draw[42][4] = 0;rain_draw[43][4] = 0;rain_draw[44][4] = 0;rain_draw[45][4] = 0;rain_draw[46][4] = 0;rain_draw[47][4] = 0;rain_draw[48][4] = 0;rain_draw[49][4] = 0;rain_draw[50][4] = 0;rain_draw[51][4] = 0;rain_draw[52][4] = 0;rain_draw[53][4] = 0;rain_draw[54][4] = 0;rain_draw[55][4] = 0;rain_draw[56][4] = 0;rain_draw[57][4] = 0;rain_draw[58][4] = 0;rain_draw[59][4] = 0;rain_draw[60][4] = 0;rain_draw[61][4] = 0;rain_draw[62][4] = 0;rain_draw[63][4] = 0;rain_draw[64][4] = 0;rain_draw[65][4] = 0;rain_draw[66][4] = 0;rain_draw[67][4] = 0;rain_draw[68][4] = 0;rain_draw[69][4] = 0;rain_draw[70][4] = 0;rain_draw[71][4] = 0;rain_draw[72][4] = 0;rain_draw[73][4] = 0;rain_draw[74][4] = 0;rain_draw[75][4] = 0;rain_draw[76][4] = 0;rain_draw[77][4] = 0;rain_draw[78][4] = 0;rain_draw[79][4] = 0;rain_draw[80][4] = 0;rain_draw[81][4] = 0;rain_draw[82][4] = 0;rain_draw[83][4] = 0;rain_draw[84][4] = 0;rain_draw[85][4] = 0;rain_draw[86][4] = 0;rain_draw[87][4] = 0;rain_draw[88][4] = 0;rain_draw[89][4] = 0;rain_draw[90][4] = 0;rain_draw[91][4] = 0;rain_draw[92][4] = 0;rain_draw[93][4] = 0;rain_draw[94][4] = 0;rain_draw[95][4] = 0;
        rain_draw[0][5] = 0;rain_draw[1][5] = 0;rain_draw[2][5] = 0;rain_draw[3][5] = 0;rain_draw[4][5] = 0;rain_draw[5][5] = 0;rain_draw[6][5] = 0;rain_draw[7][5] = 0;rain_draw[8][5] = 0;rain_draw[9][5] = 0;rain_draw[10][5] = 0;rain_draw[11][5] = 0;rain_draw[12][5] = 0;rain_draw[13][5] = 0;rain_draw[14][5] = 0;rain_draw[15][5] = 0;rain_draw[16][5] = 0;rain_draw[17][5] = 0;rain_draw[18][5] = 0;rain_draw[19][5] = 0;rain_draw[20][5] = 0;rain_draw[21][5] = 0;rain_draw[22][5] = 0;rain_draw[23][5] = 0;rain_draw[24][5] = 0;rain_draw[25][5] = 0;rain_draw[26][5] = 0;rain_draw[27][5] = 0;rain_draw[28][5] = 0;rain_draw[29][5] = 0;rain_draw[30][5] = 0;rain_draw[31][5] = 0;rain_draw[32][5] = 0;rain_draw[33][5] = 0;rain_draw[34][5] = 0;rain_draw[35][5] = 0;rain_draw[36][5] = 0;rain_draw[37][5] = 0;rain_draw[38][5] = 0;rain_draw[39][5] = 0;rain_draw[40][5] = 0;rain_draw[41][5] = 0;rain_draw[42][5] = 0;rain_draw[43][5] = 0;rain_draw[44][5] = 0;rain_draw[45][5] = 0;rain_draw[46][5] = 0;rain_draw[47][5] = 0;rain_draw[48][5] = 0;rain_draw[49][5] = 1;rain_draw[50][5] = 1;rain_draw[51][5] = 1;rain_draw[52][5] = 0;rain_draw[53][5] = 0;rain_draw[54][5] = 0;rain_draw[55][5] = 0;rain_draw[56][5] = 0;rain_draw[57][5] = 0;rain_draw[58][5] = 0;rain_draw[59][5] = 0;rain_draw[60][5] = 0;rain_draw[61][5] = 0;rain_draw[62][5] = 0;rain_draw[63][5] = 0;rain_draw[64][5] = 0;rain_draw[65][5] = 0;rain_draw[66][5] = 0;rain_draw[67][5] = 0;rain_draw[68][5] = 0;rain_draw[69][5] = 0;rain_draw[70][5] = 0;rain_draw[71][5] = 0;rain_draw[72][5] = 0;rain_draw[73][5] = 0;rain_draw[74][5] = 0;rain_draw[75][5] = 0;rain_draw[76][5] = 0;rain_draw[77][5] = 0;rain_draw[78][5] = 0;rain_draw[79][5] = 0;rain_draw[80][5] = 0;rain_draw[81][5] = 0;rain_draw[82][5] = 0;rain_draw[83][5] = 0;rain_draw[84][5] = 0;rain_draw[85][5] = 0;rain_draw[86][5] = 0;rain_draw[87][5] = 0;rain_draw[88][5] = 0;rain_draw[89][5] = 0;rain_draw[90][5] = 0;rain_draw[91][5] = 0;rain_draw[92][5] = 0;rain_draw[93][5] = 0;rain_draw[94][5] = 0;rain_draw[95][5] = 0;
        rain_draw[0][6] = 0;rain_draw[1][6] = 0;rain_draw[2][6] = 0;rain_draw[3][6] = 0;rain_draw[4][6] = 0;rain_draw[5][6] = 0;rain_draw[6][6] = 0;rain_draw[7][6] = 0;rain_draw[8][6] = 0;rain_draw[9][6] = 0;rain_draw[10][6] = 1;rain_draw[11][6] = 1;rain_draw[12][6] = 1;rain_draw[13][6] = 0;rain_draw[14][6] = 0;rain_draw[15][6] = 0;rain_draw[16][6] = 0;rain_draw[17][6] = 0;rain_draw[18][6] = 0;rain_draw[19][6] = 0;rain_draw[20][6] = 0;rain_draw[21][6] = 0;rain_draw[22][6] = 0;rain_draw[23][6] = 0;rain_draw[24][6] = 0;rain_draw[25][6] = 0;rain_draw[26][6] = 0;rain_draw[27][6] = 0;rain_draw[28][6] = 0;rain_draw[29][6] = 0;rain_draw[30][6] = 0;rain_draw[31][6] = 0;rain_draw[32][6] = 0;rain_draw[33][6] = 0;rain_draw[34][6] = 0;rain_draw[35][6] = 0;rain_draw[36][6] = 0;rain_draw[37][6] = 0;rain_draw[38][6] = 0;rain_draw[39][6] = 0;rain_draw[40][6] = 0;rain_draw[41][6] = 0;rain_draw[42][6] = 0;rain_draw[43][6] = 0;rain_draw[44][6] = 0;rain_draw[45][6] = 0;rain_draw[46][6] = 0;rain_draw[47][6] = 0;rain_draw[48][6] = 1;rain_draw[49][6] = 1;rain_draw[50][6] = 1;rain_draw[51][6] = 0;rain_draw[52][6] = 0;rain_draw[53][6] = 0;rain_draw[54][6] = 0;rain_draw[55][6] = 0;rain_draw[56][6] = 0;rain_draw[57][6] = 0;rain_draw[58][6] = 0;rain_draw[59][6] = 0;rain_draw[60][6] = 0;rain_draw[61][6] = 0;rain_draw[62][6] = 0;rain_draw[63][6] = 0;rain_draw[64][6] = 0;rain_draw[65][6] = 0;rain_draw[66][6] = 0;rain_draw[67][6] = 0;rain_draw[68][6] = 0;rain_draw[69][6] = 0;rain_draw[70][6] = 0;rain_draw[71][6] = 0;rain_draw[72][6] = 0;rain_draw[73][6] = 0;rain_draw[74][6] = 0;rain_draw[75][6] = 0;rain_draw[76][6] = 0;rain_draw[77][6] = 0;rain_draw[78][6] = 0;rain_draw[79][6] = 0;rain_draw[80][6] = 0;rain_draw[81][6] = 0;rain_draw[82][6] = 0;rain_draw[83][6] = 0;rain_draw[84][6] = 0;rain_draw[85][6] = 0;rain_draw[86][6] = 0;rain_draw[87][6] = 0;rain_draw[88][6] = 0;rain_draw[89][6] = 0;rain_draw[90][6] = 0;rain_draw[91][6] = 0;rain_draw[92][6] = 0;rain_draw[93][6] = 0;rain_draw[94][6] = 0;rain_draw[95][6] = 0;
        rain_draw[0][7] = 0;rain_draw[1][7] = 0;rain_draw[2][7] = 0;rain_draw[3][7] = 0;rain_draw[4][7] = 0;rain_draw[5][7] = 0;rain_draw[6][7] = 0;rain_draw[7][7] = 0;rain_draw[8][7] = 0;rain_draw[9][7] = 1;rain_draw[10][7] = 1;rain_draw[11][7] = 1;rain_draw[12][7] = 0;rain_draw[13][7] = 0;rain_draw[14][7] = 0;rain_draw[15][7] = 0;rain_draw[16][7] = 0;rain_draw[17][7] = 0;rain_draw[18][7] = 0;rain_draw[19][7] = 0;rain_draw[20][7] = 0;rain_draw[21][7] = 0;rain_draw[22][7] = 0;rain_draw[23][7] = 0;rain_draw[24][7] = 0;rain_draw[25][7] = 0;rain_draw[26][7] = 0;rain_draw[27][7] = 0;rain_draw[28][7] = 0;rain_draw[29][7] = 0;rain_draw[30][7] = 0;rain_draw[31][7] = 0;rain_draw[32][7] = 0;rain_draw[33][7] = 0;rain_draw[34][7] = 0;rain_draw[35][7] = 0;rain_draw[36][7] = 0;rain_draw[37][7] = 0;rain_draw[38][7] = 0;rain_draw[39][7] = 0;rain_draw[40][7] = 0;rain_draw[41][7] = 0;rain_draw[42][7] = 0;rain_draw[43][7] = 0;rain_draw[44][7] = 0;rain_draw[45][7] = 0;rain_draw[46][7] = 0;rain_draw[47][7] = 1;rain_draw[48][7] = 1;rain_draw[49][7] = 1;rain_draw[50][7] = 0;rain_draw[51][7] = 0;rain_draw[52][7] = 0;rain_draw[53][7] = 0;rain_draw[54][7] = 0;rain_draw[55][7] = 0;rain_draw[56][7] = 0;rain_draw[57][7] = 0;rain_draw[58][7] = 0;rain_draw[59][7] = 0;rain_draw[60][7] = 0;rain_draw[61][7] = 0;rain_draw[62][7] = 0;rain_draw[63][7] = 0;rain_draw[64][7] = 0;rain_draw[65][7] = 0;rain_draw[66][7] = 0;rain_draw[67][7] = 0;rain_draw[68][7] = 0;rain_draw[69][7] = 0;rain_draw[70][7] = 1;rain_draw[71][7] = 1;rain_draw[72][7] = 1;rain_draw[73][7] = 0;rain_draw[74][7] = 0;rain_draw[75][7] = 0;rain_draw[76][7] = 0;rain_draw[77][7] = 0;rain_draw[78][7] = 0;rain_draw[79][7] = 0;rain_draw[80][7] = 0;rain_draw[81][7] = 0;rain_draw[82][7] = 0;rain_draw[83][7] = 0;rain_draw[84][7] = 0;rain_draw[85][7] = 0;rain_draw[86][7] = 0;rain_draw[87][7] = 0;rain_draw[88][7] = 0;rain_draw[89][7] = 0;rain_draw[90][7] = 0;rain_draw[91][7] = 0;rain_draw[92][7] = 0;rain_draw[93][7] = 0;rain_draw[94][7] = 0;rain_draw[95][7] = 0;
        rain_draw[0][8] = 0;rain_draw[1][8] = 0;rain_draw[2][8] = 0;rain_draw[3][8] = 0;rain_draw[4][8] = 0;rain_draw[5][8] = 0;rain_draw[6][8] = 0;rain_draw[7][8] = 0;rain_draw[8][8] = 1;rain_draw[9][8] = 1;rain_draw[10][8] = 1;rain_draw[11][8] = 0;rain_draw[12][8] = 0;rain_draw[13][8] = 0;rain_draw[14][8] = 0;rain_draw[15][8] = 0;rain_draw[16][8] = 0;rain_draw[17][8] = 0;rain_draw[18][8] = 0;rain_draw[19][8] = 0;rain_draw[20][8] = 0;rain_draw[21][8] = 0;rain_draw[22][8] = 0;rain_draw[23][8] = 0;rain_draw[24][8] = 0;rain_draw[25][8] = 0;rain_draw[26][8] = 0;rain_draw[27][8] = 0;rain_draw[28][8] = 0;rain_draw[29][8] = 0;rain_draw[30][8] = 0;rain_draw[31][8] = 0;rain_draw[32][8] = 0;rain_draw[33][8] = 0;rain_draw[34][8] = 0;rain_draw[35][8] = 0;rain_draw[36][8] = 0;rain_draw[37][8] = 0;rain_draw[38][8] = 0;rain_draw[39][8] = 0;rain_draw[40][8] = 0;rain_draw[41][8] = 0;rain_draw[42][8] = 0;rain_draw[43][8] = 0;rain_draw[44][8] = 0;rain_draw[45][8] = 0;rain_draw[46][8] = 1;rain_draw[47][8] = 1;rain_draw[48][8] = 1;rain_draw[49][8] = 0;rain_draw[50][8] = 0;rain_draw[51][8] = 0;rain_draw[52][8] = 0;rain_draw[53][8] = 0;rain_draw[54][8] = 0;rain_draw[55][8] = 0;rain_draw[56][8] = 0;rain_draw[57][8] = 0;rain_draw[58][8] = 0;rain_draw[59][8] = 0;rain_draw[60][8] = 0;rain_draw[61][8] = 0;rain_draw[62][8] = 0;rain_draw[63][8] = 0;rain_draw[64][8] = 0;rain_draw[65][8] = 0;rain_draw[66][8] = 0;rain_draw[67][8] = 0;rain_draw[68][8] = 0;rain_draw[69][8] = 1;rain_draw[70][8] = 1;rain_draw[71][8] = 1;rain_draw[72][8] = 0;rain_draw[73][8] = 0;rain_draw[74][8] = 0;rain_draw[75][8] = 0;rain_draw[76][8] = 0;rain_draw[77][8] = 0;rain_draw[78][8] = 0;rain_draw[79][8] = 0;rain_draw[80][8] = 0;rain_draw[81][8] = 0;rain_draw[82][8] = 0;rain_draw[83][8] = 0;rain_draw[84][8] = 0;rain_draw[85][8] = 0;rain_draw[86][8] = 0;rain_draw[87][8] = 0;rain_draw[88][8] = 0;rain_draw[89][8] = 0;rain_draw[90][8] = 0;rain_draw[91][8] = 0;rain_draw[92][8] = 0;rain_draw[93][8] = 0;rain_draw[94][8] = 0;rain_draw[95][8] = 0;
        rain_draw[0][9] = 0;rain_draw[1][9] = 0;rain_draw[2][9] = 0;rain_draw[3][9] = 0;rain_draw[4][9] = 0;rain_draw[5][9] = 0;rain_draw[6][9] = 0;rain_draw[7][9] = 1;rain_draw[8][9] = 1;rain_draw[9][9] = 1;rain_draw[10][9] = 0;rain_draw[11][9] = 0;rain_draw[12][9] = 0;rain_draw[13][9] = 0;rain_draw[14][9] = 0;rain_draw[15][9] = 0;rain_draw[16][9] = 0;rain_draw[17][9] = 0;rain_draw[18][9] = 0;rain_draw[19][9] = 0;rain_draw[20][9] = 0;rain_draw[21][9] = 0;rain_draw[22][9] = 0;rain_draw[23][9] = 0;rain_draw[24][9] = 0;rain_draw[25][9] = 0;rain_draw[26][9] = 0;rain_draw[27][9] = 0;rain_draw[28][9] = 0;rain_draw[29][9] = 0;rain_draw[30][9] = 0;rain_draw[31][9] = 0;rain_draw[32][9] = 0;rain_draw[33][9] = 0;rain_draw[34][9] = 0;rain_draw[35][9] = 0;rain_draw[36][9] = 0;rain_draw[37][9] = 0;rain_draw[38][9] = 0;rain_draw[39][9] = 0;rain_draw[40][9] = 0;rain_draw[41][9] = 0;rain_draw[42][9] = 0;rain_draw[43][9] = 0;rain_draw[44][9] = 0;rain_draw[45][9] = 1;rain_draw[46][9] = 1;rain_draw[47][9] = 1;rain_draw[48][9] = 0;rain_draw[49][9] = 0;rain_draw[50][9] = 0;rain_draw[51][9] = 0;rain_draw[52][9] = 0;rain_draw[53][9] = 0;rain_draw[54][9] = 0;rain_draw[55][9] = 0;rain_draw[56][9] = 0;rain_draw[57][9] = 0;rain_draw[58][9] = 0;rain_draw[59][9] = 0;rain_draw[60][9] = 0;rain_draw[61][9] = 0;rain_draw[62][9] = 0;rain_draw[63][9] = 0;rain_draw[64][9] = 0;rain_draw[65][9] = 0;rain_draw[66][9] = 0;rain_draw[67][9] = 0;rain_draw[68][9] = 1;rain_draw[69][9] = 1;rain_draw[70][9] = 1;rain_draw[71][9] = 0;rain_draw[72][9] = 0;rain_draw[73][9] = 0;rain_draw[74][9] = 0;rain_draw[75][9] = 0;rain_draw[76][9] = 0;rain_draw[77][9] = 0;rain_draw[78][9] = 0;rain_draw[79][9] = 0;rain_draw[80][9] = 0;rain_draw[81][9] = 0;rain_draw[82][9] = 0;rain_draw[83][9] = 0;rain_draw[84][9] = 0;rain_draw[85][9] = 0;rain_draw[86][9] = 0;rain_draw[87][9] = 0;rain_draw[88][9] = 0;rain_draw[89][9] = 0;rain_draw[90][9] = 0;rain_draw[91][9] = 0;rain_draw[92][9] = 0;rain_draw[93][9] = 0;rain_draw[94][9] = 0;rain_draw[95][9] = 0;
        rain_draw[0][10] = 0;rain_draw[1][10] = 0;rain_draw[2][10] = 0;rain_draw[3][10] = 0;rain_draw[4][10] = 0;rain_draw[5][10] = 0;rain_draw[6][10] = 1;rain_draw[7][10] = 1;rain_draw[8][10] = 1;rain_draw[9][10] = 0;rain_draw[10][10] = 0;rain_draw[11][10] = 0;rain_draw[12][10] = 0;rain_draw[13][10] = 0;rain_draw[14][10] = 0;rain_draw[15][10] = 0;rain_draw[16][10] = 0;rain_draw[17][10] = 0;rain_draw[18][10] = 0;rain_draw[19][10] = 0;rain_draw[20][10] = 0;rain_draw[21][10] = 0;rain_draw[22][10] = 0;rain_draw[23][10] = 0;rain_draw[24][10] = 0;rain_draw[25][10] = 0;rain_draw[26][10] = 0;rain_draw[27][10] = 0;rain_draw[28][10] = 0;rain_draw[29][10] = 0;rain_draw[30][10] = 0;rain_draw[31][10] = 0;rain_draw[32][10] = 0;rain_draw[33][10] = 0;rain_draw[34][10] = 0;rain_draw[35][10] = 0;rain_draw[36][10] = 0;rain_draw[37][10] = 0;rain_draw[38][10] = 0;rain_draw[39][10] = 0;rain_draw[40][10] = 0;rain_draw[41][10] = 0;rain_draw[42][10] = 0;rain_draw[43][10] = 0;rain_draw[44][10] = 1;rain_draw[45][10] = 1;rain_draw[46][10] = 1;rain_draw[47][10] = 0;rain_draw[48][10] = 0;rain_draw[49][10] = 0;rain_draw[50][10] = 0;rain_draw[51][10] = 0;rain_draw[52][10] = 0;rain_draw[53][10] = 0;rain_draw[54][10] = 0;rain_draw[55][10] = 0;rain_draw[56][10] = 0;rain_draw[57][10] = 0;rain_draw[58][10] = 0;rain_draw[59][10] = 0;rain_draw[60][10] = 0;rain_draw[61][10] = 0;rain_draw[62][10] = 0;rain_draw[63][10] = 0;rain_draw[64][10] = 0;rain_draw[65][10] = 0;rain_draw[66][10] = 0;rain_draw[67][10] = 1;rain_draw[68][10] = 1;rain_draw[69][10] = 1;rain_draw[70][10] = 0;rain_draw[71][10] = 0;rain_draw[72][10] = 0;rain_draw[73][10] = 0;rain_draw[74][10] = 0;rain_draw[75][10] = 0;rain_draw[76][10] = 0;rain_draw[77][10] = 0;rain_draw[78][10] = 0;rain_draw[79][10] = 0;rain_draw[80][10] = 0;rain_draw[81][10] = 0;rain_draw[82][10] = 0;rain_draw[83][10] = 0;rain_draw[84][10] = 0;rain_draw[85][10] = 0;rain_draw[86][10] = 0;rain_draw[87][10] = 0;rain_draw[88][10] = 0;rain_draw[89][10] = 0;rain_draw[90][10] = 0;rain_draw[91][10] = 0;rain_draw[92][10] = 0;rain_draw[93][10] = 0;rain_draw[94][10] = 0;rain_draw[95][10] = 0;
        rain_draw[0][11] = 0;rain_draw[1][11] = 0;rain_draw[2][11] = 0;rain_draw[3][11] = 0;rain_draw[4][11] = 0;rain_draw[5][11] = 1;rain_draw[6][11] = 1;rain_draw[7][11] = 1;rain_draw[8][11] = 0;rain_draw[9][11] = 0;rain_draw[10][11] = 0;rain_draw[11][11] = 0;rain_draw[12][11] = 0;rain_draw[13][11] = 0;rain_draw[14][11] = 0;rain_draw[15][11] = 0;rain_draw[16][11] = 0;rain_draw[17][11] = 0;rain_draw[18][11] = 0;rain_draw[19][11] = 0;rain_draw[20][11] = 0;rain_draw[21][11] = 0;rain_draw[22][11] = 0;rain_draw[23][11] = 0;rain_draw[24][11] = 0;rain_draw[25][11] = 0;rain_draw[26][11] = 0;rain_draw[27][11] = 0;rain_draw[28][11] = 0;rain_draw[29][11] = 0;rain_draw[30][11] = 0;rain_draw[31][11] = 0;rain_draw[32][11] = 0;rain_draw[33][11] = 0;rain_draw[34][11] = 0;rain_draw[35][11] = 0;rain_draw[36][11] = 0;rain_draw[37][11] = 0;rain_draw[38][11] = 0;rain_draw[39][11] = 0;rain_draw[40][11] = 0;rain_draw[41][11] = 0;rain_draw[42][11] = 0;rain_draw[43][11] = 1;rain_draw[44][11] = 1;rain_draw[45][11] = 1;rain_draw[46][11] = 0;rain_draw[47][11] = 0;rain_draw[48][11] = 0;rain_draw[49][11] = 0;rain_draw[50][11] = 0;rain_draw[51][11] = 0;rain_draw[52][11] = 0;rain_draw[53][11] = 0;rain_draw[54][11] = 0;rain_draw[55][11] = 0;rain_draw[56][11] = 0;rain_draw[57][11] = 0;rain_draw[58][11] = 0;rain_draw[59][11] = 0;rain_draw[60][11] = 0;rain_draw[61][11] = 0;rain_draw[62][11] = 0;rain_draw[63][11] = 0;rain_draw[64][11] = 0;rain_draw[65][11] = 0;rain_draw[66][11] = 1;rain_draw[67][11] = 1;rain_draw[68][11] = 1;rain_draw[69][11] = 0;rain_draw[70][11] = 0;rain_draw[71][11] = 0;rain_draw[72][11] = 0;rain_draw[73][11] = 0;rain_draw[74][11] = 0;rain_draw[75][11] = 0;rain_draw[76][11] = 0;rain_draw[77][11] = 0;rain_draw[78][11] = 0;rain_draw[79][11] = 0;rain_draw[80][11] = 0;rain_draw[81][11] = 0;rain_draw[82][11] = 0;rain_draw[83][11] = 0;rain_draw[84][11] = 0;rain_draw[85][11] = 0;rain_draw[86][11] = 0;rain_draw[87][11] = 0;rain_draw[88][11] = 0;rain_draw[89][11] = 0;rain_draw[90][11] = 0;rain_draw[91][11] = 0;rain_draw[92][11] = 0;rain_draw[93][11] = 0;rain_draw[94][11] = 0;rain_draw[95][11] = 0;
        rain_draw[0][12] = 0;rain_draw[1][12] = 0;rain_draw[2][12] = 0;rain_draw[3][12] = 0;rain_draw[4][12] = 1;rain_draw[5][12] = 1;rain_draw[6][12] = 1;rain_draw[7][12] = 0;rain_draw[8][12] = 0;rain_draw[9][12] = 0;rain_draw[10][12] = 0;rain_draw[11][12] = 0;rain_draw[12][12] = 0;rain_draw[13][12] = 0;rain_draw[14][12] = 0;rain_draw[15][12] = 0;rain_draw[16][12] = 0;rain_draw[17][12] = 0;rain_draw[18][12] = 0;rain_draw[19][12] = 0;rain_draw[20][12] = 0;rain_draw[21][12] = 0;rain_draw[22][12] = 0;rain_draw[23][12] = 0;rain_draw[24][12] = 0;rain_draw[25][12] = 0;rain_draw[26][12] = 0;rain_draw[27][12] = 0;rain_draw[28][12] = 0;rain_draw[29][12] = 0;rain_draw[30][12] = 0;rain_draw[31][12] = 0;rain_draw[32][12] = 0;rain_draw[33][12] = 0;rain_draw[34][12] = 0;rain_draw[35][12] = 0;rain_draw[36][12] = 0;rain_draw[37][12] = 0;rain_draw[38][12] = 0;rain_draw[39][12] = 0;rain_draw[40][12] = 0;rain_draw[41][12] = 0;rain_draw[42][12] = 0;rain_draw[43][12] = 0;rain_draw[44][12] = 0;rain_draw[45][12] = 0;rain_draw[46][12] = 0;rain_draw[47][12] = 0;rain_draw[48][12] = 0;rain_draw[49][12] = 0;rain_draw[50][12] = 0;rain_draw[51][12] = 0;rain_draw[52][12] = 0;rain_draw[53][12] = 0;rain_draw[54][12] = 0;rain_draw[55][12] = 0;rain_draw[56][12] = 0;rain_draw[57][12] = 0;rain_draw[58][12] = 0;rain_draw[59][12] = 0;rain_draw[60][12] = 0;rain_draw[61][12] = 0;rain_draw[62][12] = 0;rain_draw[63][12] = 0;rain_draw[64][12] = 0;rain_draw[65][12] = 1;rain_draw[66][12] = 1;rain_draw[67][12] = 1;rain_draw[68][12] = 0;rain_draw[69][12] = 0;rain_draw[70][12] = 0;rain_draw[71][12] = 0;rain_draw[72][12] = 0;rain_draw[73][12] = 0;rain_draw[74][12] = 0;rain_draw[75][12] = 0;rain_draw[76][12] = 0;rain_draw[77][12] = 0;rain_draw[78][12] = 0;rain_draw[79][12] = 0;rain_draw[80][12] = 0;rain_draw[81][12] = 0;rain_draw[82][12] = 0;rain_draw[83][12] = 0;rain_draw[84][12] = 0;rain_draw[85][12] = 0;rain_draw[86][12] = 0;rain_draw[87][12] = 0;rain_draw[88][12] = 0;rain_draw[89][12] = 0;rain_draw[90][12] = 0;rain_draw[91][12] = 0;rain_draw[92][12] = 0;rain_draw[93][12] = 0;rain_draw[94][12] = 0;rain_draw[95][12] = 0;
        rain_draw[0][13] = 0;rain_draw[1][13] = 0;rain_draw[2][13] = 0;rain_draw[3][13] = 0;rain_draw[4][13] = 0;rain_draw[5][13] = 0;rain_draw[6][13] = 0;rain_draw[7][13] = 0;rain_draw[8][13] = 0;rain_draw[9][13] = 0;rain_draw[10][13] = 0;rain_draw[11][13] = 0;rain_draw[12][13] = 0;rain_draw[13][13] = 0;rain_draw[14][13] = 0;rain_draw[15][13] = 0;rain_draw[16][13] = 0;rain_draw[17][13] = 0;rain_draw[18][13] = 0;rain_draw[19][13] = 0;rain_draw[20][13] = 0;rain_draw[21][13] = 0;rain_draw[22][13] = 0;rain_draw[23][13] = 0;rain_draw[24][13] = 0;rain_draw[25][13] = 0;rain_draw[26][13] = 0;rain_draw[27][13] = 0;rain_draw[28][13] = 0;rain_draw[29][13] = 0;rain_draw[30][13] = 0;rain_draw[31][13] = 0;rain_draw[32][13] = 0;rain_draw[33][13] = 0;rain_draw[34][13] = 0;rain_draw[35][13] = 0;rain_draw[36][13] = 0;rain_draw[37][13] = 0;rain_draw[38][13] = 0;rain_draw[39][13] = 0;rain_draw[40][13] = 0;rain_draw[41][13] = 0;rain_draw[42][13] = 0;rain_draw[43][13] = 0;rain_draw[44][13] = 0;rain_draw[45][13] = 0;rain_draw[46][13] = 0;rain_draw[47][13] = 0;rain_draw[48][13] = 0;rain_draw[49][13] = 0;rain_draw[50][13] = 0;rain_draw[51][13] = 0;rain_draw[52][13] = 0;rain_draw[53][13] = 0;rain_draw[54][13] = 0;rain_draw[55][13] = 0;rain_draw[56][13] = 0;rain_draw[57][13] = 0;rain_draw[58][13] = 0;rain_draw[59][13] = 0;rain_draw[60][13] = 0;rain_draw[61][13] = 0;rain_draw[62][13] = 0;rain_draw[63][13] = 0;rain_draw[64][13] = 1;rain_draw[65][13] = 1;rain_draw[66][13] = 1;rain_draw[67][13] = 0;rain_draw[68][13] = 0;rain_draw[69][13] = 0;rain_draw[70][13] = 0;rain_draw[71][13] = 0;rain_draw[72][13] = 0;rain_draw[73][13] = 0;rain_draw[74][13] = 0;rain_draw[75][13] = 0;rain_draw[76][13] = 0;rain_draw[77][13] = 0;rain_draw[78][13] = 0;rain_draw[79][13] = 0;rain_draw[80][13] = 0;rain_draw[81][13] = 0;rain_draw[82][13] = 0;rain_draw[83][13] = 0;rain_draw[84][13] = 0;rain_draw[85][13] = 0;rain_draw[86][13] = 0;rain_draw[87][13] = 0;rain_draw[88][13] = 0;rain_draw[89][13] = 0;rain_draw[90][13] = 0;rain_draw[91][13] = 0;rain_draw[92][13] = 0;rain_draw[93][13] = 0;rain_draw[94][13] = 0;rain_draw[95][13] = 0;
        rain_draw[0][14] = 0;rain_draw[1][14] = 0;rain_draw[2][14] = 0;rain_draw[3][14] = 0;rain_draw[4][14] = 0;rain_draw[5][14] = 0;rain_draw[6][14] = 0;rain_draw[7][14] = 0;rain_draw[8][14] = 0;rain_draw[9][14] = 0;rain_draw[10][14] = 0;rain_draw[11][14] = 0;rain_draw[12][14] = 0;rain_draw[13][14] = 0;rain_draw[14][14] = 0;rain_draw[15][14] = 0;rain_draw[16][14] = 0;rain_draw[17][14] = 0;rain_draw[18][14] = 0;rain_draw[19][14] = 0;rain_draw[20][14] = 0;rain_draw[21][14] = 0;rain_draw[22][14] = 0;rain_draw[23][14] = 0;rain_draw[24][14] = 0;rain_draw[25][14] = 0;rain_draw[26][14] = 0;rain_draw[27][14] = 0;rain_draw[28][14] = 0;rain_draw[29][14] = 0;rain_draw[30][14] = 0;rain_draw[31][14] = 0;rain_draw[32][14] = 0;rain_draw[33][14] = 0;rain_draw[34][14] = 0;rain_draw[35][14] = 0;rain_draw[36][14] = 0;rain_draw[37][14] = 0;rain_draw[38][14] = 0;rain_draw[39][14] = 0;rain_draw[40][14] = 0;rain_draw[41][14] = 0;rain_draw[42][14] = 0;rain_draw[43][14] = 0;rain_draw[44][14] = 0;rain_draw[45][14] = 0;rain_draw[46][14] = 0;rain_draw[47][14] = 0;rain_draw[48][14] = 0;rain_draw[49][14] = 0;rain_draw[50][14] = 0;rain_draw[51][14] = 0;rain_draw[52][14] = 0;rain_draw[53][14] = 0;rain_draw[54][14] = 0;rain_draw[55][14] = 0;rain_draw[56][14] = 0;rain_draw[57][14] = 0;rain_draw[58][14] = 0;rain_draw[59][14] = 0;rain_draw[60][14] = 0;rain_draw[61][14] = 0;rain_draw[62][14] = 0;rain_draw[63][14] = 0;rain_draw[64][14] = 0;rain_draw[65][14] = 0;rain_draw[66][14] = 0;rain_draw[67][14] = 0;rain_draw[68][14] = 0;rain_draw[69][14] = 0;rain_draw[70][14] = 0;rain_draw[71][14] = 0;rain_draw[72][14] = 0;rain_draw[73][14] = 0;rain_draw[74][14] = 0;rain_draw[75][14] = 0;rain_draw[76][14] = 0;rain_draw[77][14] = 0;rain_draw[78][14] = 0;rain_draw[79][14] = 0;rain_draw[80][14] = 0;rain_draw[81][14] = 0;rain_draw[82][14] = 0;rain_draw[83][14] = 0;rain_draw[84][14] = 1;rain_draw[85][14] = 1;rain_draw[86][14] = 1;rain_draw[87][14] = 0;rain_draw[88][14] = 0;rain_draw[89][14] = 0;rain_draw[90][14] = 0;rain_draw[91][14] = 0;rain_draw[92][14] = 0;rain_draw[93][14] = 0;rain_draw[94][14] = 0;rain_draw[95][14] = 0;
        rain_draw[0][15] = 0;rain_draw[1][15] = 0;rain_draw[2][15] = 0;rain_draw[3][15] = 0;rain_draw[4][15] = 0;rain_draw[5][15] = 0;rain_draw[6][15] = 0;rain_draw[7][15] = 0;rain_draw[8][15] = 0;rain_draw[9][15] = 0;rain_draw[10][15] = 0;rain_draw[11][15] = 0;rain_draw[12][15] = 0;rain_draw[13][15] = 0;rain_draw[14][15] = 0;rain_draw[15][15] = 0;rain_draw[16][15] = 0;rain_draw[17][15] = 0;rain_draw[18][15] = 0;rain_draw[19][15] = 0;rain_draw[20][15] = 0;rain_draw[21][15] = 0;rain_draw[22][15] = 0;rain_draw[23][15] = 0;rain_draw[24][15] = 0;rain_draw[25][15] = 0;rain_draw[26][15] = 0;rain_draw[27][15] = 0;rain_draw[28][15] = 0;rain_draw[29][15] = 0;rain_draw[30][15] = 0;rain_draw[31][15] = 0;rain_draw[32][15] = 0;rain_draw[33][15] = 0;rain_draw[34][15] = 0;rain_draw[35][15] = 0;rain_draw[36][15] = 0;rain_draw[37][15] = 0;rain_draw[38][15] = 0;rain_draw[39][15] = 0;rain_draw[40][15] = 0;rain_draw[41][15] = 0;rain_draw[42][15] = 0;rain_draw[43][15] = 0;rain_draw[44][15] = 0;rain_draw[45][15] = 0;rain_draw[46][15] = 0;rain_draw[47][15] = 0;rain_draw[48][15] = 0;rain_draw[49][15] = 0;rain_draw[50][15] = 0;rain_draw[51][15] = 0;rain_draw[52][15] = 0;rain_draw[53][15] = 0;rain_draw[54][15] = 0;rain_draw[55][15] = 0;rain_draw[56][15] = 0;rain_draw[57][15] = 0;rain_draw[58][15] = 0;rain_draw[59][15] = 0;rain_draw[60][15] = 0;rain_draw[61][15] = 0;rain_draw[62][15] = 0;rain_draw[63][15] = 0;rain_draw[64][15] = 0;rain_draw[65][15] = 0;rain_draw[66][15] = 0;rain_draw[67][15] = 0;rain_draw[68][15] = 0;rain_draw[69][15] = 0;rain_draw[70][15] = 0;rain_draw[71][15] = 0;rain_draw[72][15] = 0;rain_draw[73][15] = 0;rain_draw[74][15] = 0;rain_draw[75][15] = 0;rain_draw[76][15] = 0;rain_draw[77][15] = 0;rain_draw[78][15] = 0;rain_draw[79][15] = 0;rain_draw[80][15] = 0;rain_draw[81][15] = 0;rain_draw[82][15] = 0;rain_draw[83][15] = 1;rain_draw[84][15] = 1;rain_draw[85][15] = 1;rain_draw[86][15] = 0;rain_draw[87][15] = 0;rain_draw[88][15] = 0;rain_draw[89][15] = 0;rain_draw[90][15] = 0;rain_draw[91][15] = 0;rain_draw[92][15] = 0;rain_draw[93][15] = 0;rain_draw[94][15] = 0;rain_draw[95][15] = 0;
        rain_draw[0][16] = 0;rain_draw[1][16] = 0;rain_draw[2][16] = 0;rain_draw[3][16] = 0;rain_draw[4][16] = 0;rain_draw[5][16] = 0;rain_draw[6][16] = 0;rain_draw[7][16] = 0;rain_draw[8][16] = 0;rain_draw[9][16] = 0;rain_draw[10][16] = 0;rain_draw[11][16] = 0;rain_draw[12][16] = 0;rain_draw[13][16] = 0;rain_draw[14][16] = 0;rain_draw[15][16] = 0;rain_draw[16][16] = 0;rain_draw[17][16] = 0;rain_draw[18][16] = 0;rain_draw[19][16] = 0;rain_draw[20][16] = 0;rain_draw[21][16] = 0;rain_draw[22][16] = 0;rain_draw[23][16] = 0;rain_draw[24][16] = 0;rain_draw[25][16] = 0;rain_draw[26][16] = 0;rain_draw[27][16] = 0;rain_draw[28][16] = 0;rain_draw[29][16] = 0;rain_draw[30][16] = 0;rain_draw[31][16] = 0;rain_draw[32][16] = 0;rain_draw[33][16] = 0;rain_draw[34][16] = 0;rain_draw[35][16] = 0;rain_draw[36][16] = 0;rain_draw[37][16] = 0;rain_draw[38][16] = 0;rain_draw[39][16] = 0;rain_draw[40][16] = 0;rain_draw[41][16] = 0;rain_draw[42][16] = 0;rain_draw[43][16] = 0;rain_draw[44][16] = 0;rain_draw[45][16] = 0;rain_draw[46][16] = 0;rain_draw[47][16] = 0;rain_draw[48][16] = 0;rain_draw[49][16] = 0;rain_draw[50][16] = 0;rain_draw[51][16] = 0;rain_draw[52][16] = 0;rain_draw[53][16] = 0;rain_draw[54][16] = 0;rain_draw[55][16] = 0;rain_draw[56][16] = 0;rain_draw[57][16] = 0;rain_draw[58][16] = 0;rain_draw[59][16] = 0;rain_draw[60][16] = 0;rain_draw[61][16] = 0;rain_draw[62][16] = 0;rain_draw[63][16] = 0;rain_draw[64][16] = 0;rain_draw[65][16] = 0;rain_draw[66][16] = 0;rain_draw[67][16] = 0;rain_draw[68][16] = 0;rain_draw[69][16] = 0;rain_draw[70][16] = 0;rain_draw[71][16] = 0;rain_draw[72][16] = 0;rain_draw[73][16] = 0;rain_draw[74][16] = 0;rain_draw[75][16] = 0;rain_draw[76][16] = 0;rain_draw[77][16] = 0;rain_draw[78][16] = 0;rain_draw[79][16] = 0;rain_draw[80][16] = 0;rain_draw[81][16] = 0;rain_draw[82][16] = 1;rain_draw[83][16] = 1;rain_draw[84][16] = 1;rain_draw[85][16] = 0;rain_draw[86][16] = 0;rain_draw[87][16] = 0;rain_draw[88][16] = 0;rain_draw[89][16] = 0;rain_draw[90][16] = 0;rain_draw[91][16] = 0;rain_draw[92][16] = 0;rain_draw[93][16] = 0;rain_draw[94][16] = 0;rain_draw[95][16] = 0;
        rain_draw[0][17] = 0;rain_draw[1][17] = 0;rain_draw[2][17] = 0;rain_draw[3][17] = 0;rain_draw[4][17] = 0;rain_draw[5][17] = 0;rain_draw[6][17] = 0;rain_draw[7][17] = 0;rain_draw[8][17] = 0;rain_draw[9][17] = 0;rain_draw[10][17] = 0;rain_draw[11][17] = 0;rain_draw[12][17] = 0;rain_draw[13][17] = 0;rain_draw[14][17] = 0;rain_draw[15][17] = 0;rain_draw[16][17] = 0;rain_draw[17][17] = 0;rain_draw[18][17] = 0;rain_draw[19][17] = 0;rain_draw[20][17] = 0;rain_draw[21][17] = 0;rain_draw[22][17] = 0;rain_draw[23][17] = 0;rain_draw[24][17] = 0;rain_draw[25][17] = 0;rain_draw[26][17] = 0;rain_draw[27][17] = 0;rain_draw[28][17] = 0;rain_draw[29][17] = 0;rain_draw[30][17] = 0;rain_draw[31][17] = 0;rain_draw[32][17] = 0;rain_draw[33][17] = 0;rain_draw[34][17] = 0;rain_draw[35][17] = 0;rain_draw[36][17] = 0;rain_draw[37][17] = 0;rain_draw[38][17] = 0;rain_draw[39][17] = 0;rain_draw[40][17] = 0;rain_draw[41][17] = 0;rain_draw[42][17] = 0;rain_draw[43][17] = 0;rain_draw[44][17] = 0;rain_draw[45][17] = 0;rain_draw[46][17] = 0;rain_draw[47][17] = 0;rain_draw[48][17] = 0;rain_draw[49][17] = 0;rain_draw[50][17] = 0;rain_draw[51][17] = 0;rain_draw[52][17] = 0;rain_draw[53][17] = 0;rain_draw[54][17] = 0;rain_draw[55][17] = 0;rain_draw[56][17] = 0;rain_draw[57][17] = 0;rain_draw[58][17] = 0;rain_draw[59][17] = 0;rain_draw[60][17] = 0;rain_draw[61][17] = 0;rain_draw[62][17] = 0;rain_draw[63][17] = 0;rain_draw[64][17] = 0;rain_draw[65][17] = 0;rain_draw[66][17] = 0;rain_draw[67][17] = 0;rain_draw[68][17] = 0;rain_draw[69][17] = 0;rain_draw[70][17] = 0;rain_draw[71][17] = 0;rain_draw[72][17] = 0;rain_draw[73][17] = 0;rain_draw[74][17] = 0;rain_draw[75][17] = 0;rain_draw[76][17] = 0;rain_draw[77][17] = 0;rain_draw[78][17] = 0;rain_draw[79][17] = 0;rain_draw[80][17] = 0;rain_draw[81][17] = 1;rain_draw[82][17] = 1;rain_draw[83][17] = 1;rain_draw[84][17] = 0;rain_draw[85][17] = 0;rain_draw[86][17] = 0;rain_draw[87][17] = 0;rain_draw[88][17] = 0;rain_draw[89][17] = 0;rain_draw[90][17] = 0;rain_draw[91][17] = 0;rain_draw[92][17] = 0;rain_draw[93][17] = 0;rain_draw[94][17] = 0;rain_draw[95][17] = 0;
        rain_draw[0][18] = 0;rain_draw[1][18] = 0;rain_draw[2][18] = 0;rain_draw[3][18] = 0;rain_draw[4][18] = 0;rain_draw[5][18] = 0;rain_draw[6][18] = 0;rain_draw[7][18] = 0;rain_draw[8][18] = 0;rain_draw[9][18] = 0;rain_draw[10][18] = 0;rain_draw[11][18] = 0;rain_draw[12][18] = 0;rain_draw[13][18] = 0;rain_draw[14][18] = 0;rain_draw[15][18] = 0;rain_draw[16][18] = 0;rain_draw[17][18] = 0;rain_draw[18][18] = 0;rain_draw[19][18] = 0;rain_draw[20][18] = 0;rain_draw[21][18] = 0;rain_draw[22][18] = 0;rain_draw[23][18] = 0;rain_draw[24][18] = 0;rain_draw[25][18] = 0;rain_draw[26][18] = 0;rain_draw[27][18] = 0;rain_draw[28][18] = 1;rain_draw[29][18] = 1;rain_draw[30][18] = 1;rain_draw[31][18] = 0;rain_draw[32][18] = 0;rain_draw[33][18] = 0;rain_draw[34][18] = 0;rain_draw[35][18] = 0;rain_draw[36][18] = 0;rain_draw[37][18] = 0;rain_draw[38][18] = 0;rain_draw[39][18] = 0;rain_draw[40][18] = 0;rain_draw[41][18] = 0;rain_draw[42][18] = 0;rain_draw[43][18] = 0;rain_draw[44][18] = 0;rain_draw[45][18] = 0;rain_draw[46][18] = 0;rain_draw[47][18] = 0;rain_draw[48][18] = 0;rain_draw[49][18] = 0;rain_draw[50][18] = 0;rain_draw[51][18] = 0;rain_draw[52][18] = 0;rain_draw[53][18] = 0;rain_draw[54][18] = 0;rain_draw[55][18] = 0;rain_draw[56][18] = 0;rain_draw[57][18] = 0;rain_draw[58][18] = 0;rain_draw[59][18] = 0;rain_draw[60][18] = 0;rain_draw[61][18] = 0;rain_draw[62][18] = 0;rain_draw[63][18] = 0;rain_draw[64][18] = 0;rain_draw[65][18] = 0;rain_draw[66][18] = 0;rain_draw[67][18] = 0;rain_draw[68][18] = 0;rain_draw[69][18] = 0;rain_draw[70][18] = 0;rain_draw[71][18] = 0;rain_draw[72][18] = 0;rain_draw[73][18] = 0;rain_draw[74][18] = 0;rain_draw[75][18] = 0;rain_draw[76][18] = 0;rain_draw[77][18] = 0;rain_draw[78][18] = 0;rain_draw[79][18] = 0;rain_draw[80][18] = 1;rain_draw[81][18] = 1;rain_draw[82][18] = 1;rain_draw[83][18] = 0;rain_draw[84][18] = 0;rain_draw[85][18] = 0;rain_draw[86][18] = 0;rain_draw[87][18] = 0;rain_draw[88][18] = 0;rain_draw[89][18] = 0;rain_draw[90][18] = 0;rain_draw[91][18] = 0;rain_draw[92][18] = 0;rain_draw[93][18] = 0;rain_draw[94][18] = 0;rain_draw[95][18] = 0;
        rain_draw[0][19] = 0;rain_draw[1][19] = 0;rain_draw[2][19] = 0;rain_draw[3][19] = 0;rain_draw[4][19] = 0;rain_draw[5][19] = 0;rain_draw[6][19] = 0;rain_draw[7][19] = 0;rain_draw[8][19] = 0;rain_draw[9][19] = 0;rain_draw[10][19] = 0;rain_draw[11][19] = 0;rain_draw[12][19] = 0;rain_draw[13][19] = 0;rain_draw[14][19] = 0;rain_draw[15][19] = 0;rain_draw[16][19] = 0;rain_draw[17][19] = 0;rain_draw[18][19] = 0;rain_draw[19][19] = 0;rain_draw[20][19] = 0;rain_draw[21][19] = 0;rain_draw[22][19] = 0;rain_draw[23][19] = 0;rain_draw[24][19] = 0;rain_draw[25][19] = 0;rain_draw[26][19] = 0;rain_draw[27][19] = 1;rain_draw[28][19] = 1;rain_draw[29][19] = 1;rain_draw[30][19] = 0;rain_draw[31][19] = 0;rain_draw[32][19] = 0;rain_draw[33][19] = 0;rain_draw[34][19] = 0;rain_draw[35][19] = 0;rain_draw[36][19] = 0;rain_draw[37][19] = 0;rain_draw[38][19] = 0;rain_draw[39][19] = 0;rain_draw[40][19] = 0;rain_draw[41][19] = 0;rain_draw[42][19] = 0;rain_draw[43][19] = 0;rain_draw[44][19] = 0;rain_draw[45][19] = 0;rain_draw[46][19] = 0;rain_draw[47][19] = 0;rain_draw[48][19] = 0;rain_draw[49][19] = 0;rain_draw[50][19] = 0;rain_draw[51][19] = 0;rain_draw[52][19] = 0;rain_draw[53][19] = 0;rain_draw[54][19] = 0;rain_draw[55][19] = 0;rain_draw[56][19] = 0;rain_draw[57][19] = 0;rain_draw[58][19] = 0;rain_draw[59][19] = 0;rain_draw[60][19] = 0;rain_draw[61][19] = 0;rain_draw[62][19] = 0;rain_draw[63][19] = 0;rain_draw[64][19] = 0;rain_draw[65][19] = 0;rain_draw[66][19] = 0;rain_draw[67][19] = 0;rain_draw[68][19] = 0;rain_draw[69][19] = 0;rain_draw[70][19] = 0;rain_draw[71][19] = 0;rain_draw[72][19] = 0;rain_draw[73][19] = 0;rain_draw[74][19] = 0;rain_draw[75][19] = 0;rain_draw[76][19] = 0;rain_draw[77][19] = 0;rain_draw[78][19] = 0;rain_draw[79][19] = 1;rain_draw[80][19] = 1;rain_draw[81][19] = 1;rain_draw[82][19] = 0;rain_draw[83][19] = 0;rain_draw[84][19] = 0;rain_draw[85][19] = 0;rain_draw[86][19] = 0;rain_draw[87][19] = 0;rain_draw[88][19] = 0;rain_draw[89][19] = 0;rain_draw[90][19] = 0;rain_draw[91][19] = 0;rain_draw[92][19] = 0;rain_draw[93][19] = 0;rain_draw[94][19] = 0;rain_draw[95][19] = 0;
        rain_draw[0][20] = 0;rain_draw[1][20] = 0;rain_draw[2][20] = 0;rain_draw[3][20] = 0;rain_draw[4][20] = 0;rain_draw[5][20] = 0;rain_draw[6][20] = 0;rain_draw[7][20] = 0;rain_draw[8][20] = 0;rain_draw[9][20] = 0;rain_draw[10][20] = 0;rain_draw[11][20] = 0;rain_draw[12][20] = 0;rain_draw[13][20] = 0;rain_draw[14][20] = 0;rain_draw[15][20] = 0;rain_draw[16][20] = 0;rain_draw[17][20] = 0;rain_draw[18][20] = 0;rain_draw[19][20] = 0;rain_draw[20][20] = 0;rain_draw[21][20] = 0;rain_draw[22][20] = 0;rain_draw[23][20] = 0;rain_draw[24][20] = 0;rain_draw[25][20] = 0;rain_draw[26][20] = 1;rain_draw[27][20] = 1;rain_draw[28][20] = 1;rain_draw[29][20] = 0;rain_draw[30][20] = 0;rain_draw[31][20] = 0;rain_draw[32][20] = 0;rain_draw[33][20] = 0;rain_draw[34][20] = 0;rain_draw[35][20] = 0;rain_draw[36][20] = 0;rain_draw[37][20] = 0;rain_draw[38][20] = 0;rain_draw[39][20] = 0;rain_draw[40][20] = 0;rain_draw[41][20] = 0;rain_draw[42][20] = 0;rain_draw[43][20] = 0;rain_draw[44][20] = 0;rain_draw[45][20] = 0;rain_draw[46][20] = 0;rain_draw[47][20] = 0;rain_draw[48][20] = 0;rain_draw[49][20] = 0;rain_draw[50][20] = 0;rain_draw[51][20] = 0;rain_draw[52][20] = 0;rain_draw[53][20] = 0;rain_draw[54][20] = 0;rain_draw[55][20] = 0;rain_draw[56][20] = 0;rain_draw[57][20] = 0;rain_draw[58][20] = 0;rain_draw[59][20] = 0;rain_draw[60][20] = 0;rain_draw[61][20] = 0;rain_draw[62][20] = 0;rain_draw[63][20] = 0;rain_draw[64][20] = 0;rain_draw[65][20] = 0;rain_draw[66][20] = 0;rain_draw[67][20] = 0;rain_draw[68][20] = 0;rain_draw[69][20] = 0;rain_draw[70][20] = 0;rain_draw[71][20] = 0;rain_draw[72][20] = 0;rain_draw[73][20] = 0;rain_draw[74][20] = 0;rain_draw[75][20] = 0;rain_draw[76][20] = 0;rain_draw[77][20] = 0;rain_draw[78][20] = 1;rain_draw[79][20] = 1;rain_draw[80][20] = 1;rain_draw[81][20] = 0;rain_draw[82][20] = 0;rain_draw[83][20] = 0;rain_draw[84][20] = 0;rain_draw[85][20] = 0;rain_draw[86][20] = 0;rain_draw[87][20] = 0;rain_draw[88][20] = 0;rain_draw[89][20] = 0;rain_draw[90][20] = 0;rain_draw[91][20] = 0;rain_draw[92][20] = 0;rain_draw[93][20] = 0;rain_draw[94][20] = 0;rain_draw[95][20] = 0;
        rain_draw[0][21] = 0;rain_draw[1][21] = 0;rain_draw[2][21] = 0;rain_draw[3][21] = 0;rain_draw[4][21] = 0;rain_draw[5][21] = 0;rain_draw[6][21] = 0;rain_draw[7][21] = 0;rain_draw[8][21] = 0;rain_draw[9][21] = 0;rain_draw[10][21] = 0;rain_draw[11][21] = 0;rain_draw[12][21] = 0;rain_draw[13][21] = 0;rain_draw[14][21] = 0;rain_draw[15][21] = 0;rain_draw[16][21] = 0;rain_draw[17][21] = 0;rain_draw[18][21] = 0;rain_draw[19][21] = 0;rain_draw[20][21] = 0;rain_draw[21][21] = 0;rain_draw[22][21] = 0;rain_draw[23][21] = 0;rain_draw[24][21] = 0;rain_draw[25][21] = 1;rain_draw[26][21] = 1;rain_draw[27][21] = 1;rain_draw[28][21] = 0;rain_draw[29][21] = 0;rain_draw[30][21] = 0;rain_draw[31][21] = 0;rain_draw[32][21] = 0;rain_draw[33][21] = 0;rain_draw[34][21] = 0;rain_draw[35][21] = 0;rain_draw[36][21] = 0;rain_draw[37][21] = 0;rain_draw[38][21] = 0;rain_draw[39][21] = 0;rain_draw[40][21] = 0;rain_draw[41][21] = 0;rain_draw[42][21] = 0;rain_draw[43][21] = 0;rain_draw[44][21] = 0;rain_draw[45][21] = 0;rain_draw[46][21] = 0;rain_draw[47][21] = 0;rain_draw[48][21] = 0;rain_draw[49][21] = 0;rain_draw[50][21] = 0;rain_draw[51][21] = 0;rain_draw[52][21] = 0;rain_draw[53][21] = 0;rain_draw[54][21] = 0;rain_draw[55][21] = 0;rain_draw[56][21] = 0;rain_draw[57][21] = 0;rain_draw[58][21] = 0;rain_draw[59][21] = 0;rain_draw[60][21] = 0;rain_draw[61][21] = 0;rain_draw[62][21] = 0;rain_draw[63][21] = 0;rain_draw[64][21] = 0;rain_draw[65][21] = 0;rain_draw[66][21] = 0;rain_draw[67][21] = 0;rain_draw[68][21] = 0;rain_draw[69][21] = 0;rain_draw[70][21] = 0;rain_draw[71][21] = 0;rain_draw[72][21] = 0;rain_draw[73][21] = 0;rain_draw[74][21] = 0;rain_draw[75][21] = 0;rain_draw[76][21] = 0;rain_draw[77][21] = 0;rain_draw[78][21] = 0;rain_draw[79][21] = 0;rain_draw[80][21] = 0;rain_draw[81][21] = 0;rain_draw[82][21] = 0;rain_draw[83][21] = 0;rain_draw[84][21] = 0;rain_draw[85][21] = 0;rain_draw[86][21] = 0;rain_draw[87][21] = 0;rain_draw[88][21] = 0;rain_draw[89][21] = 0;rain_draw[90][21] = 0;rain_draw[91][21] = 0;rain_draw[92][21] = 0;rain_draw[93][21] = 0;rain_draw[94][21] = 0;rain_draw[95][21] = 0;
        rain_draw[0][22] = 0;rain_draw[1][22] = 0;rain_draw[2][22] = 0;rain_draw[3][22] = 0;rain_draw[4][22] = 0;rain_draw[5][22] = 0;rain_draw[6][22] = 0;rain_draw[7][22] = 0;rain_draw[8][22] = 0;rain_draw[9][22] = 0;rain_draw[10][22] = 0;rain_draw[11][22] = 0;rain_draw[12][22] = 0;rain_draw[13][22] = 0;rain_draw[14][22] = 0;rain_draw[15][22] = 0;rain_draw[16][22] = 0;rain_draw[17][22] = 0;rain_draw[18][22] = 0;rain_draw[19][22] = 0;rain_draw[20][22] = 0;rain_draw[21][22] = 0;rain_draw[22][22] = 0;rain_draw[23][22] = 0;rain_draw[24][22] = 1;rain_draw[25][22] = 1;rain_draw[26][22] = 1;rain_draw[27][22] = 0;rain_draw[28][22] = 0;rain_draw[29][22] = 0;rain_draw[30][22] = 0;rain_draw[31][22] = 0;rain_draw[32][22] = 0;rain_draw[33][22] = 0;rain_draw[34][22] = 0;rain_draw[35][22] = 0;rain_draw[36][22] = 0;rain_draw[37][22] = 0;rain_draw[38][22] = 0;rain_draw[39][22] = 0;rain_draw[40][22] = 0;rain_draw[41][22] = 0;rain_draw[42][22] = 0;rain_draw[43][22] = 0;rain_draw[44][22] = 0;rain_draw[45][22] = 0;rain_draw[46][22] = 0;rain_draw[47][22] = 0;rain_draw[48][22] = 0;rain_draw[49][22] = 0;rain_draw[50][22] = 0;rain_draw[51][22] = 0;rain_draw[52][22] = 0;rain_draw[53][22] = 0;rain_draw[54][22] = 0;rain_draw[55][22] = 0;rain_draw[56][22] = 0;rain_draw[57][22] = 0;rain_draw[58][22] = 0;rain_draw[59][22] = 0;rain_draw[60][22] = 0;rain_draw[61][22] = 0;rain_draw[62][22] = 0;rain_draw[63][22] = 0;rain_draw[64][22] = 0;rain_draw[65][22] = 0;rain_draw[66][22] = 0;rain_draw[67][22] = 0;rain_draw[68][22] = 0;rain_draw[69][22] = 0;rain_draw[70][22] = 0;rain_draw[71][22] = 0;rain_draw[72][22] = 0;rain_draw[73][22] = 0;rain_draw[74][22] = 0;rain_draw[75][22] = 0;rain_draw[76][22] = 0;rain_draw[77][22] = 0;rain_draw[78][22] = 0;rain_draw[79][22] = 0;rain_draw[80][22] = 0;rain_draw[81][22] = 0;rain_draw[82][22] = 0;rain_draw[83][22] = 0;rain_draw[84][22] = 0;rain_draw[85][22] = 0;rain_draw[86][22] = 0;rain_draw[87][22] = 0;rain_draw[88][22] = 0;rain_draw[89][22] = 0;rain_draw[90][22] = 0;rain_draw[91][22] = 0;rain_draw[92][22] = 0;rain_draw[93][22] = 0;rain_draw[94][22] = 0;rain_draw[95][22] = 0;
        rain_draw[0][23] = 0;rain_draw[1][23] = 0;rain_draw[2][23] = 0;rain_draw[3][23] = 0;rain_draw[4][23] = 0;rain_draw[5][23] = 0;rain_draw[6][23] = 0;rain_draw[7][23] = 0;rain_draw[8][23] = 0;rain_draw[9][23] = 0;rain_draw[10][23] = 0;rain_draw[11][23] = 0;rain_draw[12][23] = 0;rain_draw[13][23] = 0;rain_draw[14][23] = 0;rain_draw[15][23] = 0;rain_draw[16][23] = 0;rain_draw[17][23] = 0;rain_draw[18][23] = 0;rain_draw[19][23] = 0;rain_draw[20][23] = 0;rain_draw[21][23] = 0;rain_draw[22][23] = 0;rain_draw[23][23] = 1;rain_draw[24][23] = 1;rain_draw[25][23] = 1;rain_draw[26][23] = 0;rain_draw[27][23] = 0;rain_draw[28][23] = 0;rain_draw[29][23] = 0;rain_draw[30][23] = 0;rain_draw[31][23] = 0;rain_draw[32][23] = 0;rain_draw[33][23] = 0;rain_draw[34][23] = 0;rain_draw[35][23] = 0;rain_draw[36][23] = 0;rain_draw[37][23] = 0;rain_draw[38][23] = 0;rain_draw[39][23] = 0;rain_draw[40][23] = 0;rain_draw[41][23] = 0;rain_draw[42][23] = 0;rain_draw[43][23] = 0;rain_draw[44][23] = 0;rain_draw[45][23] = 0;rain_draw[46][23] = 0;rain_draw[47][23] = 0;rain_draw[48][23] = 0;rain_draw[49][23] = 0;rain_draw[50][23] = 0;rain_draw[51][23] = 0;rain_draw[52][23] = 0;rain_draw[53][23] = 0;rain_draw[54][23] = 0;rain_draw[55][23] = 0;rain_draw[56][23] = 0;rain_draw[57][23] = 0;rain_draw[58][23] = 0;rain_draw[59][23] = 0;rain_draw[60][23] = 0;rain_draw[61][23] = 0;rain_draw[62][23] = 0;rain_draw[63][23] = 0;rain_draw[64][23] = 0;rain_draw[65][23] = 0;rain_draw[66][23] = 0;rain_draw[67][23] = 0;rain_draw[68][23] = 0;rain_draw[69][23] = 0;rain_draw[70][23] = 0;rain_draw[71][23] = 0;rain_draw[72][23] = 0;rain_draw[73][23] = 0;rain_draw[74][23] = 0;rain_draw[75][23] = 0;rain_draw[76][23] = 0;rain_draw[77][23] = 0;rain_draw[78][23] = 0;rain_draw[79][23] = 0;rain_draw[80][23] = 0;rain_draw[81][23] = 0;rain_draw[82][23] = 0;rain_draw[83][23] = 0;rain_draw[84][23] = 0;rain_draw[85][23] = 0;rain_draw[86][23] = 0;rain_draw[87][23] = 0;rain_draw[88][23] = 0;rain_draw[89][23] = 0;rain_draw[90][23] = 0;rain_draw[91][23] = 0;rain_draw[92][23] = 0;rain_draw[93][23] = 0;rain_draw[94][23] = 0;rain_draw[95][23] = 0;
        rain_draw[0][24] = 0;rain_draw[1][24] = 0;rain_draw[2][24] = 0;rain_draw[3][24] = 0;rain_draw[4][24] = 0;rain_draw[5][24] = 0;rain_draw[6][24] = 0;rain_draw[7][24] = 0;rain_draw[8][24] = 0;rain_draw[9][24] = 0;rain_draw[10][24] = 0;rain_draw[11][24] = 0;rain_draw[12][24] = 0;rain_draw[13][24] = 0;rain_draw[14][24] = 0;rain_draw[15][24] = 0;rain_draw[16][24] = 0;rain_draw[17][24] = 0;rain_draw[18][24] = 0;rain_draw[19][24] = 0;rain_draw[20][24] = 0;rain_draw[21][24] = 0;rain_draw[22][24] = 1;rain_draw[23][24] = 1;rain_draw[24][24] = 1;rain_draw[25][24] = 0;rain_draw[26][24] = 0;rain_draw[27][24] = 0;rain_draw[28][24] = 0;rain_draw[29][24] = 0;rain_draw[30][24] = 0;rain_draw[31][24] = 0;rain_draw[32][24] = 0;rain_draw[33][24] = 0;rain_draw[34][24] = 0;rain_draw[35][24] = 0;rain_draw[36][24] = 0;rain_draw[37][24] = 0;rain_draw[38][24] = 0;rain_draw[39][24] = 0;rain_draw[40][24] = 0;rain_draw[41][24] = 0;rain_draw[42][24] = 0;rain_draw[43][24] = 0;rain_draw[44][24] = 0;rain_draw[45][24] = 0;rain_draw[46][24] = 0;rain_draw[47][24] = 0;rain_draw[48][24] = 0;rain_draw[49][24] = 0;rain_draw[50][24] = 0;rain_draw[51][24] = 0;rain_draw[52][24] = 0;rain_draw[53][24] = 0;rain_draw[54][24] = 0;rain_draw[55][24] = 0;rain_draw[56][24] = 0;rain_draw[57][24] = 0;rain_draw[58][24] = 0;rain_draw[59][24] = 0;rain_draw[60][24] = 0;rain_draw[61][24] = 0;rain_draw[62][24] = 0;rain_draw[63][24] = 1;rain_draw[64][24] = 1;rain_draw[65][24] = 1;rain_draw[66][24] = 0;rain_draw[67][24] = 0;rain_draw[68][24] = 0;rain_draw[69][24] = 0;rain_draw[70][24] = 0;rain_draw[71][24] = 0;rain_draw[72][24] = 0;rain_draw[73][24] = 0;rain_draw[74][24] = 0;rain_draw[75][24] = 0;rain_draw[76][24] = 0;rain_draw[77][24] = 0;rain_draw[78][24] = 0;rain_draw[79][24] = 0;rain_draw[80][24] = 0;rain_draw[81][24] = 0;rain_draw[82][24] = 0;rain_draw[83][24] = 0;rain_draw[84][24] = 0;rain_draw[85][24] = 0;rain_draw[86][24] = 0;rain_draw[87][24] = 0;rain_draw[88][24] = 0;rain_draw[89][24] = 0;rain_draw[90][24] = 0;rain_draw[91][24] = 0;rain_draw[92][24] = 0;rain_draw[93][24] = 0;rain_draw[94][24] = 0;rain_draw[95][24] = 0;
        rain_draw[0][25] = 0;rain_draw[1][25] = 0;rain_draw[2][25] = 0;rain_draw[3][25] = 0;rain_draw[4][25] = 0;rain_draw[5][25] = 0;rain_draw[6][25] = 0;rain_draw[7][25] = 0;rain_draw[8][25] = 0;rain_draw[9][25] = 0;rain_draw[10][25] = 0;rain_draw[11][25] = 0;rain_draw[12][25] = 0;rain_draw[13][25] = 0;rain_draw[14][25] = 0;rain_draw[15][25] = 0;rain_draw[16][25] = 0;rain_draw[17][25] = 0;rain_draw[18][25] = 0;rain_draw[19][25] = 0;rain_draw[20][25] = 0;rain_draw[21][25] = 0;rain_draw[22][25] = 0;rain_draw[23][25] = 0;rain_draw[24][25] = 0;rain_draw[25][25] = 0;rain_draw[26][25] = 0;rain_draw[27][25] = 0;rain_draw[28][25] = 0;rain_draw[29][25] = 0;rain_draw[30][25] = 0;rain_draw[31][25] = 0;rain_draw[32][25] = 0;rain_draw[33][25] = 0;rain_draw[34][25] = 0;rain_draw[35][25] = 0;rain_draw[36][25] = 0;rain_draw[37][25] = 0;rain_draw[38][25] = 0;rain_draw[39][25] = 0;rain_draw[40][25] = 0;rain_draw[41][25] = 0;rain_draw[42][25] = 0;rain_draw[43][25] = 0;rain_draw[44][25] = 0;rain_draw[45][25] = 1;rain_draw[46][25] = 1;rain_draw[47][25] = 1;rain_draw[48][25] = 0;rain_draw[49][25] = 0;rain_draw[50][25] = 0;rain_draw[51][25] = 0;rain_draw[52][25] = 0;rain_draw[53][25] = 0;rain_draw[54][25] = 0;rain_draw[55][25] = 0;rain_draw[56][25] = 0;rain_draw[57][25] = 0;rain_draw[58][25] = 0;rain_draw[59][25] = 0;rain_draw[60][25] = 0;rain_draw[61][25] = 0;rain_draw[62][25] = 1;rain_draw[63][25] = 1;rain_draw[64][25] = 1;rain_draw[65][25] = 0;rain_draw[66][25] = 0;rain_draw[67][25] = 0;rain_draw[68][25] = 0;rain_draw[69][25] = 0;rain_draw[70][25] = 0;rain_draw[71][25] = 0;rain_draw[72][25] = 0;rain_draw[73][25] = 0;rain_draw[74][25] = 0;rain_draw[75][25] = 0;rain_draw[76][25] = 0;rain_draw[77][25] = 0;rain_draw[78][25] = 0;rain_draw[79][25] = 0;rain_draw[80][25] = 0;rain_draw[81][25] = 0;rain_draw[82][25] = 0;rain_draw[83][25] = 0;rain_draw[84][25] = 0;rain_draw[85][25] = 0;rain_draw[86][25] = 0;rain_draw[87][25] = 0;rain_draw[88][25] = 0;rain_draw[89][25] = 0;rain_draw[90][25] = 0;rain_draw[91][25] = 0;rain_draw[92][25] = 0;rain_draw[93][25] = 0;rain_draw[94][25] = 0;rain_draw[95][25] = 0;
        rain_draw[0][26] = 0;rain_draw[1][26] = 0;rain_draw[2][26] = 0;rain_draw[3][26] = 0;rain_draw[4][26] = 0;rain_draw[5][26] = 0;rain_draw[6][26] = 0;rain_draw[7][26] = 0;rain_draw[8][26] = 0;rain_draw[9][26] = 0;rain_draw[10][26] = 0;rain_draw[11][26] = 0;rain_draw[12][26] = 0;rain_draw[13][26] = 0;rain_draw[14][26] = 0;rain_draw[15][26] = 0;rain_draw[16][26] = 0;rain_draw[17][26] = 0;rain_draw[18][26] = 0;rain_draw[19][26] = 0;rain_draw[20][26] = 0;rain_draw[21][26] = 0;rain_draw[22][26] = 0;rain_draw[23][26] = 0;rain_draw[24][26] = 0;rain_draw[25][26] = 0;rain_draw[26][26] = 0;rain_draw[27][26] = 0;rain_draw[28][26] = 0;rain_draw[29][26] = 0;rain_draw[30][26] = 0;rain_draw[31][26] = 0;rain_draw[32][26] = 0;rain_draw[33][26] = 0;rain_draw[34][26] = 0;rain_draw[35][26] = 0;rain_draw[36][26] = 0;rain_draw[37][26] = 0;rain_draw[38][26] = 0;rain_draw[39][26] = 0;rain_draw[40][26] = 0;rain_draw[41][26] = 0;rain_draw[42][26] = 0;rain_draw[43][26] = 0;rain_draw[44][26] = 1;rain_draw[45][26] = 1;rain_draw[46][26] = 1;rain_draw[47][26] = 0;rain_draw[48][26] = 0;rain_draw[49][26] = 0;rain_draw[50][26] = 0;rain_draw[51][26] = 0;rain_draw[52][26] = 0;rain_draw[53][26] = 0;rain_draw[54][26] = 0;rain_draw[55][26] = 0;rain_draw[56][26] = 0;rain_draw[57][26] = 0;rain_draw[58][26] = 0;rain_draw[59][26] = 0;rain_draw[60][26] = 0;rain_draw[61][26] = 1;rain_draw[62][26] = 1;rain_draw[63][26] = 1;rain_draw[64][26] = 0;rain_draw[65][26] = 0;rain_draw[66][26] = 0;rain_draw[67][26] = 0;rain_draw[68][26] = 0;rain_draw[69][26] = 0;rain_draw[70][26] = 0;rain_draw[71][26] = 0;rain_draw[72][26] = 0;rain_draw[73][26] = 0;rain_draw[74][26] = 0;rain_draw[75][26] = 0;rain_draw[76][26] = 0;rain_draw[77][26] = 0;rain_draw[78][26] = 0;rain_draw[79][26] = 0;rain_draw[80][26] = 0;rain_draw[81][26] = 0;rain_draw[82][26] = 0;rain_draw[83][26] = 0;rain_draw[84][26] = 0;rain_draw[85][26] = 0;rain_draw[86][26] = 0;rain_draw[87][26] = 0;rain_draw[88][26] = 0;rain_draw[89][26] = 0;rain_draw[90][26] = 0;rain_draw[91][26] = 0;rain_draw[92][26] = 0;rain_draw[93][26] = 0;rain_draw[94][26] = 0;rain_draw[95][26] = 0;
        rain_draw[0][27] = 0;rain_draw[1][27] = 0;rain_draw[2][27] = 0;rain_draw[3][27] = 0;rain_draw[4][27] = 0;rain_draw[5][27] = 0;rain_draw[6][27] = 0;rain_draw[7][27] = 0;rain_draw[8][27] = 0;rain_draw[9][27] = 0;rain_draw[10][27] = 0;rain_draw[11][27] = 0;rain_draw[12][27] = 0;rain_draw[13][27] = 0;rain_draw[14][27] = 0;rain_draw[15][27] = 0;rain_draw[16][27] = 0;rain_draw[17][27] = 0;rain_draw[18][27] = 0;rain_draw[19][27] = 0;rain_draw[20][27] = 0;rain_draw[21][27] = 0;rain_draw[22][27] = 0;rain_draw[23][27] = 0;rain_draw[24][27] = 0;rain_draw[25][27] = 0;rain_draw[26][27] = 0;rain_draw[27][27] = 0;rain_draw[28][27] = 0;rain_draw[29][27] = 0;rain_draw[30][27] = 0;rain_draw[31][27] = 0;rain_draw[32][27] = 0;rain_draw[33][27] = 0;rain_draw[34][27] = 0;rain_draw[35][27] = 0;rain_draw[36][27] = 0;rain_draw[37][27] = 0;rain_draw[38][27] = 0;rain_draw[39][27] = 0;rain_draw[40][27] = 0;rain_draw[41][27] = 0;rain_draw[42][27] = 0;rain_draw[43][27] = 1;rain_draw[44][27] = 1;rain_draw[45][27] = 1;rain_draw[46][27] = 0;rain_draw[47][27] = 0;rain_draw[48][27] = 0;rain_draw[49][27] = 0;rain_draw[50][27] = 0;rain_draw[51][27] = 0;rain_draw[52][27] = 0;rain_draw[53][27] = 0;rain_draw[54][27] = 0;rain_draw[55][27] = 0;rain_draw[56][27] = 0;rain_draw[57][27] = 0;rain_draw[58][27] = 0;rain_draw[59][27] = 0;rain_draw[60][27] = 1;rain_draw[61][27] = 1;rain_draw[62][27] = 1;rain_draw[63][27] = 0;rain_draw[64][27] = 0;rain_draw[65][27] = 0;rain_draw[66][27] = 0;rain_draw[67][27] = 0;rain_draw[68][27] = 0;rain_draw[69][27] = 0;rain_draw[70][27] = 0;rain_draw[71][27] = 0;rain_draw[72][27] = 0;rain_draw[73][27] = 0;rain_draw[74][27] = 0;rain_draw[75][27] = 0;rain_draw[76][27] = 0;rain_draw[77][27] = 0;rain_draw[78][27] = 0;rain_draw[79][27] = 0;rain_draw[80][27] = 0;rain_draw[81][27] = 0;rain_draw[82][27] = 0;rain_draw[83][27] = 0;rain_draw[84][27] = 0;rain_draw[85][27] = 0;rain_draw[86][27] = 0;rain_draw[87][27] = 0;rain_draw[88][27] = 0;rain_draw[89][27] = 0;rain_draw[90][27] = 0;rain_draw[91][27] = 0;rain_draw[92][27] = 0;rain_draw[93][27] = 0;rain_draw[94][27] = 0;rain_draw[95][27] = 0;
        rain_draw[0][28] = 0;rain_draw[1][28] = 0;rain_draw[2][28] = 0;rain_draw[3][28] = 0;rain_draw[4][28] = 0;rain_draw[5][28] = 0;rain_draw[6][28] = 0;rain_draw[7][28] = 0;rain_draw[8][28] = 0;rain_draw[9][28] = 0;rain_draw[10][28] = 0;rain_draw[11][28] = 0;rain_draw[12][28] = 0;rain_draw[13][28] = 0;rain_draw[14][28] = 0;rain_draw[15][28] = 0;rain_draw[16][28] = 0;rain_draw[17][28] = 0;rain_draw[18][28] = 0;rain_draw[19][28] = 0;rain_draw[20][28] = 0;rain_draw[21][28] = 0;rain_draw[22][28] = 0;rain_draw[23][28] = 0;rain_draw[24][28] = 0;rain_draw[25][28] = 0;rain_draw[26][28] = 0;rain_draw[27][28] = 0;rain_draw[28][28] = 0;rain_draw[29][28] = 0;rain_draw[30][28] = 0;rain_draw[31][28] = 0;rain_draw[32][28] = 0;rain_draw[33][28] = 0;rain_draw[34][28] = 0;rain_draw[35][28] = 0;rain_draw[36][28] = 0;rain_draw[37][28] = 0;rain_draw[38][28] = 0;rain_draw[39][28] = 0;rain_draw[40][28] = 0;rain_draw[41][28] = 0;rain_draw[42][28] = 1;rain_draw[43][28] = 1;rain_draw[44][28] = 1;rain_draw[45][28] = 0;rain_draw[46][28] = 0;rain_draw[47][28] = 0;rain_draw[48][28] = 0;rain_draw[49][28] = 0;rain_draw[50][28] = 0;rain_draw[51][28] = 0;rain_draw[52][28] = 0;rain_draw[53][28] = 0;rain_draw[54][28] = 0;rain_draw[55][28] = 0;rain_draw[56][28] = 0;rain_draw[57][28] = 0;rain_draw[58][28] = 0;rain_draw[59][28] = 1;rain_draw[60][28] = 1;rain_draw[61][28] = 1;rain_draw[62][28] = 0;rain_draw[63][28] = 0;rain_draw[64][28] = 0;rain_draw[65][28] = 0;rain_draw[66][28] = 0;rain_draw[67][28] = 0;rain_draw[68][28] = 0;rain_draw[69][28] = 0;rain_draw[70][28] = 0;rain_draw[71][28] = 0;rain_draw[72][28] = 0;rain_draw[73][28] = 0;rain_draw[74][28] = 0;rain_draw[75][28] = 0;rain_draw[76][28] = 0;rain_draw[77][28] = 0;rain_draw[78][28] = 0;rain_draw[79][28] = 0;rain_draw[80][28] = 0;rain_draw[81][28] = 0;rain_draw[82][28] = 0;rain_draw[83][28] = 0;rain_draw[84][28] = 0;rain_draw[85][28] = 0;rain_draw[86][28] = 0;rain_draw[87][28] = 0;rain_draw[88][28] = 0;rain_draw[89][28] = 0;rain_draw[90][28] = 0;rain_draw[91][28] = 0;rain_draw[92][28] = 0;rain_draw[93][28] = 0;rain_draw[94][28] = 0;rain_draw[95][28] = 0;
        rain_draw[0][29] = 0;rain_draw[1][29] = 0;rain_draw[2][29] = 0;rain_draw[3][29] = 0;rain_draw[4][29] = 0;rain_draw[5][29] = 0;rain_draw[6][29] = 0;rain_draw[7][29] = 0;rain_draw[8][29] = 0;rain_draw[9][29] = 0;rain_draw[10][29] = 0;rain_draw[11][29] = 1;rain_draw[12][29] = 1;rain_draw[13][29] = 1;rain_draw[14][29] = 0;rain_draw[15][29] = 0;rain_draw[16][29] = 0;rain_draw[17][29] = 0;rain_draw[18][29] = 0;rain_draw[19][29] = 0;rain_draw[20][29] = 0;rain_draw[21][29] = 0;rain_draw[22][29] = 0;rain_draw[23][29] = 0;rain_draw[24][29] = 0;rain_draw[25][29] = 0;rain_draw[26][29] = 0;rain_draw[27][29] = 0;rain_draw[28][29] = 0;rain_draw[29][29] = 0;rain_draw[30][29] = 0;rain_draw[31][29] = 0;rain_draw[32][29] = 0;rain_draw[33][29] = 0;rain_draw[34][29] = 0;rain_draw[35][29] = 0;rain_draw[36][29] = 0;rain_draw[37][29] = 0;rain_draw[38][29] = 0;rain_draw[39][29] = 0;rain_draw[40][29] = 0;rain_draw[41][29] = 1;rain_draw[42][29] = 1;rain_draw[43][29] = 1;rain_draw[44][29] = 0;rain_draw[45][29] = 0;rain_draw[46][29] = 0;rain_draw[47][29] = 0;rain_draw[48][29] = 0;rain_draw[49][29] = 0;rain_draw[50][29] = 0;rain_draw[51][29] = 0;rain_draw[52][29] = 0;rain_draw[53][29] = 0;rain_draw[54][29] = 0;rain_draw[55][29] = 0;rain_draw[56][29] = 0;rain_draw[57][29] = 0;rain_draw[58][29] = 1;rain_draw[59][29] = 1;rain_draw[60][29] = 1;rain_draw[61][29] = 0;rain_draw[62][29] = 0;rain_draw[63][29] = 0;rain_draw[64][29] = 0;rain_draw[65][29] = 0;rain_draw[66][29] = 0;rain_draw[67][29] = 0;rain_draw[68][29] = 0;rain_draw[69][29] = 0;rain_draw[70][29] = 0;rain_draw[71][29] = 0;rain_draw[72][29] = 0;rain_draw[73][29] = 0;rain_draw[74][29] = 0;rain_draw[75][29] = 0;rain_draw[76][29] = 0;rain_draw[77][29] = 0;rain_draw[78][29] = 0;rain_draw[79][29] = 0;rain_draw[80][29] = 0;rain_draw[81][29] = 0;rain_draw[82][29] = 0;rain_draw[83][29] = 0;rain_draw[84][29] = 0;rain_draw[85][29] = 0;rain_draw[86][29] = 0;rain_draw[87][29] = 0;rain_draw[88][29] = 0;rain_draw[89][29] = 0;rain_draw[90][29] = 0;rain_draw[91][29] = 0;rain_draw[92][29] = 0;rain_draw[93][29] = 0;rain_draw[94][29] = 0;rain_draw[95][29] = 0;
        rain_draw[0][30] = 0;rain_draw[1][30] = 0;rain_draw[2][30] = 0;rain_draw[3][30] = 0;rain_draw[4][30] = 0;rain_draw[5][30] = 0;rain_draw[6][30] = 0;rain_draw[7][30] = 0;rain_draw[8][30] = 0;rain_draw[9][30] = 0;rain_draw[10][30] = 1;rain_draw[11][30] = 1;rain_draw[12][30] = 1;rain_draw[13][30] = 0;rain_draw[14][30] = 0;rain_draw[15][30] = 0;rain_draw[16][30] = 0;rain_draw[17][30] = 0;rain_draw[18][30] = 0;rain_draw[19][30] = 0;rain_draw[20][30] = 0;rain_draw[21][30] = 0;rain_draw[22][30] = 0;rain_draw[23][30] = 0;rain_draw[24][30] = 0;rain_draw[25][30] = 0;rain_draw[26][30] = 0;rain_draw[27][30] = 0;rain_draw[28][30] = 0;rain_draw[29][30] = 0;rain_draw[30][30] = 0;rain_draw[31][30] = 0;rain_draw[32][30] = 0;rain_draw[33][30] = 0;rain_draw[34][30] = 0;rain_draw[35][30] = 0;rain_draw[36][30] = 0;rain_draw[37][30] = 0;rain_draw[38][30] = 0;rain_draw[39][30] = 0;rain_draw[40][30] = 1;rain_draw[41][30] = 1;rain_draw[42][30] = 1;rain_draw[43][30] = 0;rain_draw[44][30] = 0;rain_draw[45][30] = 0;rain_draw[46][30] = 0;rain_draw[47][30] = 0;rain_draw[48][30] = 0;rain_draw[49][30] = 0;rain_draw[50][30] = 0;rain_draw[51][30] = 0;rain_draw[52][30] = 0;rain_draw[53][30] = 0;rain_draw[54][30] = 0;rain_draw[55][30] = 0;rain_draw[56][30] = 0;rain_draw[57][30] = 1;rain_draw[58][30] = 1;rain_draw[59][30] = 1;rain_draw[60][30] = 0;rain_draw[61][30] = 0;rain_draw[62][30] = 0;rain_draw[63][30] = 0;rain_draw[64][30] = 0;rain_draw[65][30] = 0;rain_draw[66][30] = 0;rain_draw[67][30] = 0;rain_draw[68][30] = 0;rain_draw[69][30] = 0;rain_draw[70][30] = 0;rain_draw[71][30] = 0;rain_draw[72][30] = 0;rain_draw[73][30] = 0;rain_draw[74][30] = 0;rain_draw[75][30] = 0;rain_draw[76][30] = 0;rain_draw[77][30] = 0;rain_draw[78][30] = 0;rain_draw[79][30] = 0;rain_draw[80][30] = 0;rain_draw[81][30] = 0;rain_draw[82][30] = 0;rain_draw[83][30] = 0;rain_draw[84][30] = 0;rain_draw[85][30] = 0;rain_draw[86][30] = 0;rain_draw[87][30] = 0;rain_draw[88][30] = 0;rain_draw[89][30] = 0;rain_draw[90][30] = 0;rain_draw[91][30] = 0;rain_draw[92][30] = 0;rain_draw[93][30] = 0;rain_draw[94][30] = 0;rain_draw[95][30] = 0;
        rain_draw[0][31] = 0;rain_draw[1][31] = 0;rain_draw[2][31] = 0;rain_draw[3][31] = 0;rain_draw[4][31] = 0;rain_draw[5][31] = 0;rain_draw[6][31] = 0;rain_draw[7][31] = 0;rain_draw[8][31] = 0;rain_draw[9][31] = 1;rain_draw[10][31] = 1;rain_draw[11][31] = 1;rain_draw[12][31] = 0;rain_draw[13][31] = 0;rain_draw[14][31] = 0;rain_draw[15][31] = 0;rain_draw[16][31] = 0;rain_draw[17][31] = 0;rain_draw[18][31] = 0;rain_draw[19][31] = 0;rain_draw[20][31] = 0;rain_draw[21][31] = 0;rain_draw[22][31] = 0;rain_draw[23][31] = 0;rain_draw[24][31] = 0;rain_draw[25][31] = 0;rain_draw[26][31] = 0;rain_draw[27][31] = 0;rain_draw[28][31] = 0;rain_draw[29][31] = 0;rain_draw[30][31] = 0;rain_draw[31][31] = 0;rain_draw[32][31] = 0;rain_draw[33][31] = 0;rain_draw[34][31] = 0;rain_draw[35][31] = 0;rain_draw[36][31] = 0;rain_draw[37][31] = 0;rain_draw[38][31] = 0;rain_draw[39][31] = 1;rain_draw[40][31] = 1;rain_draw[41][31] = 1;rain_draw[42][31] = 0;rain_draw[43][31] = 0;rain_draw[44][31] = 0;rain_draw[45][31] = 0;rain_draw[46][31] = 0;rain_draw[47][31] = 0;rain_draw[48][31] = 0;rain_draw[49][31] = 0;rain_draw[50][31] = 0;rain_draw[51][31] = 0;rain_draw[52][31] = 0;rain_draw[53][31] = 0;rain_draw[54][31] = 0;rain_draw[55][31] = 0;rain_draw[56][31] = 0;rain_draw[57][31] = 0;rain_draw[58][31] = 0;rain_draw[59][31] = 0;rain_draw[60][31] = 0;rain_draw[61][31] = 0;rain_draw[62][31] = 0;rain_draw[63][31] = 0;rain_draw[64][31] = 0;rain_draw[65][31] = 0;rain_draw[66][31] = 0;rain_draw[67][31] = 0;rain_draw[68][31] = 0;rain_draw[69][31] = 0;rain_draw[70][31] = 0;rain_draw[71][31] = 0;rain_draw[72][31] = 0;rain_draw[73][31] = 0;rain_draw[74][31] = 0;rain_draw[75][31] = 0;rain_draw[76][31] = 0;rain_draw[77][31] = 0;rain_draw[78][31] = 0;rain_draw[79][31] = 0;rain_draw[80][31] = 0;rain_draw[81][31] = 0;rain_draw[82][31] = 0;rain_draw[83][31] = 0;rain_draw[84][31] = 0;rain_draw[85][31] = 0;rain_draw[86][31] = 0;rain_draw[87][31] = 0;rain_draw[88][31] = 0;rain_draw[89][31] = 0;rain_draw[90][31] = 0;rain_draw[91][31] = 0;rain_draw[92][31] = 0;rain_draw[93][31] = 0;rain_draw[94][31] = 0;rain_draw[95][31] = 0;
        rain_draw[0][32] = 0;rain_draw[1][32] = 0;rain_draw[2][32] = 0;rain_draw[3][32] = 0;rain_draw[4][32] = 0;rain_draw[5][32] = 0;rain_draw[6][32] = 0;rain_draw[7][32] = 0;rain_draw[8][32] = 1;rain_draw[9][32] = 1;rain_draw[10][32] = 1;rain_draw[11][32] = 0;rain_draw[12][32] = 0;rain_draw[13][32] = 0;rain_draw[14][32] = 0;rain_draw[15][32] = 0;rain_draw[16][32] = 0;rain_draw[17][32] = 0;rain_draw[18][32] = 0;rain_draw[19][32] = 0;rain_draw[20][32] = 0;rain_draw[21][32] = 0;rain_draw[22][32] = 0;rain_draw[23][32] = 0;rain_draw[24][32] = 0;rain_draw[25][32] = 0;rain_draw[26][32] = 0;rain_draw[27][32] = 0;rain_draw[28][32] = 0;rain_draw[29][32] = 0;rain_draw[30][32] = 0;rain_draw[31][32] = 0;rain_draw[32][32] = 0;rain_draw[33][32] = 0;rain_draw[34][32] = 0;rain_draw[35][32] = 0;rain_draw[36][32] = 0;rain_draw[37][32] = 0;rain_draw[38][32] = 0;rain_draw[39][32] = 0;rain_draw[40][32] = 0;rain_draw[41][32] = 0;rain_draw[42][32] = 0;rain_draw[43][32] = 0;rain_draw[44][32] = 0;rain_draw[45][32] = 0;rain_draw[46][32] = 0;rain_draw[47][32] = 0;rain_draw[48][32] = 0;rain_draw[49][32] = 0;rain_draw[50][32] = 0;rain_draw[51][32] = 0;rain_draw[52][32] = 0;rain_draw[53][32] = 0;rain_draw[54][32] = 0;rain_draw[55][32] = 0;rain_draw[56][32] = 0;rain_draw[57][32] = 0;rain_draw[58][32] = 0;rain_draw[59][32] = 0;rain_draw[60][32] = 0;rain_draw[61][32] = 0;rain_draw[62][32] = 0;rain_draw[63][32] = 0;rain_draw[64][32] = 0;rain_draw[65][32] = 0;rain_draw[66][32] = 0;rain_draw[67][32] = 0;rain_draw[68][32] = 0;rain_draw[69][32] = 0;rain_draw[70][32] = 0;rain_draw[71][32] = 0;rain_draw[72][32] = 0;rain_draw[73][32] = 0;rain_draw[74][32] = 0;rain_draw[75][32] = 0;rain_draw[76][32] = 0;rain_draw[77][32] = 0;rain_draw[78][32] = 0;rain_draw[79][32] = 0;rain_draw[80][32] = 0;rain_draw[81][32] = 0;rain_draw[82][32] = 0;rain_draw[83][32] = 0;rain_draw[84][32] = 0;rain_draw[85][32] = 0;rain_draw[86][32] = 0;rain_draw[87][32] = 0;rain_draw[88][32] = 0;rain_draw[89][32] = 0;rain_draw[90][32] = 0;rain_draw[91][32] = 0;rain_draw[92][32] = 0;rain_draw[93][32] = 0;rain_draw[94][32] = 0;rain_draw[95][32] = 0;
        rain_draw[0][33] = 0;rain_draw[1][33] = 0;rain_draw[2][33] = 0;rain_draw[3][33] = 0;rain_draw[4][33] = 0;rain_draw[5][33] = 0;rain_draw[6][33] = 0;rain_draw[7][33] = 1;rain_draw[8][33] = 1;rain_draw[9][33] = 1;rain_draw[10][33] = 0;rain_draw[11][33] = 0;rain_draw[12][33] = 0;rain_draw[13][33] = 0;rain_draw[14][33] = 0;rain_draw[15][33] = 0;rain_draw[16][33] = 0;rain_draw[17][33] = 0;rain_draw[18][33] = 0;rain_draw[19][33] = 0;rain_draw[20][33] = 0;rain_draw[21][33] = 0;rain_draw[22][33] = 0;rain_draw[23][33] = 0;rain_draw[24][33] = 0;rain_draw[25][33] = 0;rain_draw[26][33] = 0;rain_draw[27][33] = 0;rain_draw[28][33] = 0;rain_draw[29][33] = 0;rain_draw[30][33] = 0;rain_draw[31][33] = 0;rain_draw[32][33] = 0;rain_draw[33][33] = 0;rain_draw[34][33] = 0;rain_draw[35][33] = 0;rain_draw[36][33] = 0;rain_draw[37][33] = 0;rain_draw[38][33] = 0;rain_draw[39][33] = 0;rain_draw[40][33] = 0;rain_draw[41][33] = 0;rain_draw[42][33] = 0;rain_draw[43][33] = 0;rain_draw[44][33] = 0;rain_draw[45][33] = 0;rain_draw[46][33] = 0;rain_draw[47][33] = 0;rain_draw[48][33] = 0;rain_draw[49][33] = 0;rain_draw[50][33] = 0;rain_draw[51][33] = 0;rain_draw[52][33] = 0;rain_draw[53][33] = 0;rain_draw[54][33] = 0;rain_draw[55][33] = 0;rain_draw[56][33] = 0;rain_draw[57][33] = 0;rain_draw[58][33] = 0;rain_draw[59][33] = 0;rain_draw[60][33] = 0;rain_draw[61][33] = 0;rain_draw[62][33] = 0;rain_draw[63][33] = 0;rain_draw[64][33] = 0;rain_draw[65][33] = 0;rain_draw[66][33] = 0;rain_draw[67][33] = 0;rain_draw[68][33] = 0;rain_draw[69][33] = 0;rain_draw[70][33] = 0;rain_draw[71][33] = 0;rain_draw[72][33] = 0;rain_draw[73][33] = 0;rain_draw[74][33] = 0;rain_draw[75][33] = 0;rain_draw[76][33] = 0;rain_draw[77][33] = 0;rain_draw[78][33] = 0;rain_draw[79][33] = 0;rain_draw[80][33] = 0;rain_draw[81][33] = 0;rain_draw[82][33] = 0;rain_draw[83][33] = 0;rain_draw[84][33] = 0;rain_draw[85][33] = 0;rain_draw[86][33] = 0;rain_draw[87][33] = 0;rain_draw[88][33] = 0;rain_draw[89][33] = 0;rain_draw[90][33] = 0;rain_draw[91][33] = 0;rain_draw[92][33] = 0;rain_draw[93][33] = 0;rain_draw[94][33] = 0;rain_draw[95][33] = 0;
        rain_draw[0][34] = 0;rain_draw[1][34] = 0;rain_draw[2][34] = 0;rain_draw[3][34] = 0;rain_draw[4][34] = 0;rain_draw[5][34] = 0;rain_draw[6][34] = 1;rain_draw[7][34] = 1;rain_draw[8][34] = 1;rain_draw[9][34] = 0;rain_draw[10][34] = 0;rain_draw[11][34] = 0;rain_draw[12][34] = 0;rain_draw[13][34] = 0;rain_draw[14][34] = 0;rain_draw[15][34] = 0;rain_draw[16][34] = 0;rain_draw[17][34] = 0;rain_draw[18][34] = 0;rain_draw[19][34] = 0;rain_draw[20][34] = 0;rain_draw[21][34] = 0;rain_draw[22][34] = 0;rain_draw[23][34] = 0;rain_draw[24][34] = 0;rain_draw[25][34] = 0;rain_draw[26][34] = 0;rain_draw[27][34] = 0;rain_draw[28][34] = 0;rain_draw[29][34] = 0;rain_draw[30][34] = 0;rain_draw[31][34] = 0;rain_draw[32][34] = 0;rain_draw[33][34] = 0;rain_draw[34][34] = 0;rain_draw[35][34] = 0;rain_draw[36][34] = 0;rain_draw[37][34] = 0;rain_draw[38][34] = 0;rain_draw[39][34] = 0;rain_draw[40][34] = 0;rain_draw[41][34] = 0;rain_draw[42][34] = 0;rain_draw[43][34] = 0;rain_draw[44][34] = 0;rain_draw[45][34] = 0;rain_draw[46][34] = 0;rain_draw[47][34] = 0;rain_draw[48][34] = 0;rain_draw[49][34] = 0;rain_draw[50][34] = 0;rain_draw[51][34] = 0;rain_draw[52][34] = 0;rain_draw[53][34] = 0;rain_draw[54][34] = 0;rain_draw[55][34] = 0;rain_draw[56][34] = 0;rain_draw[57][34] = 0;rain_draw[58][34] = 0;rain_draw[59][34] = 0;rain_draw[60][34] = 0;rain_draw[61][34] = 0;rain_draw[62][34] = 0;rain_draw[63][34] = 0;rain_draw[64][34] = 0;rain_draw[65][34] = 0;rain_draw[66][34] = 0;rain_draw[67][34] = 0;rain_draw[68][34] = 0;rain_draw[69][34] = 0;rain_draw[70][34] = 0;rain_draw[71][34] = 0;rain_draw[72][34] = 0;rain_draw[73][34] = 0;rain_draw[74][34] = 0;rain_draw[75][34] = 0;rain_draw[76][34] = 0;rain_draw[77][34] = 0;rain_draw[78][34] = 0;rain_draw[79][34] = 0;rain_draw[80][34] = 0;rain_draw[81][34] = 0;rain_draw[82][34] = 0;rain_draw[83][34] = 0;rain_draw[84][34] = 0;rain_draw[85][34] = 0;rain_draw[86][34] = 0;rain_draw[87][34] = 0;rain_draw[88][34] = 0;rain_draw[89][34] = 0;rain_draw[90][34] = 0;rain_draw[91][34] = 0;rain_draw[92][34] = 0;rain_draw[93][34] = 0;rain_draw[94][34] = 0;rain_draw[95][34] = 0;
        rain_draw[0][35] = 0;rain_draw[1][35] = 0;rain_draw[2][35] = 0;rain_draw[3][35] = 0;rain_draw[4][35] = 0;rain_draw[5][35] = 1;rain_draw[6][35] = 1;rain_draw[7][35] = 1;rain_draw[8][35] = 0;rain_draw[9][35] = 0;rain_draw[10][35] = 0;rain_draw[11][35] = 0;rain_draw[12][35] = 0;rain_draw[13][35] = 0;rain_draw[14][35] = 0;rain_draw[15][35] = 0;rain_draw[16][35] = 0;rain_draw[17][35] = 0;rain_draw[18][35] = 0;rain_draw[19][35] = 0;rain_draw[20][35] = 0;rain_draw[21][35] = 0;rain_draw[22][35] = 0;rain_draw[23][35] = 0;rain_draw[24][35] = 0;rain_draw[25][35] = 0;rain_draw[26][35] = 0;rain_draw[27][35] = 0;rain_draw[28][35] = 0;rain_draw[29][35] = 0;rain_draw[30][35] = 0;rain_draw[31][35] = 0;rain_draw[32][35] = 0;rain_draw[33][35] = 0;rain_draw[34][35] = 0;rain_draw[35][35] = 0;rain_draw[36][35] = 0;rain_draw[37][35] = 0;rain_draw[38][35] = 0;rain_draw[39][35] = 0;rain_draw[40][35] = 0;rain_draw[41][35] = 0;rain_draw[42][35] = 0;rain_draw[43][35] = 0;rain_draw[44][35] = 0;rain_draw[45][35] = 0;rain_draw[46][35] = 0;rain_draw[47][35] = 0;rain_draw[48][35] = 0;rain_draw[49][35] = 0;rain_draw[50][35] = 0;rain_draw[51][35] = 0;rain_draw[52][35] = 0;rain_draw[53][35] = 0;rain_draw[54][35] = 0;rain_draw[55][35] = 0;rain_draw[56][35] = 0;rain_draw[57][35] = 0;rain_draw[58][35] = 0;rain_draw[59][35] = 0;rain_draw[60][35] = 0;rain_draw[61][35] = 0;rain_draw[62][35] = 0;rain_draw[63][35] = 0;rain_draw[64][35] = 0;rain_draw[65][35] = 0;rain_draw[66][35] = 0;rain_draw[67][35] = 0;rain_draw[68][35] = 0;rain_draw[69][35] = 0;rain_draw[70][35] = 0;rain_draw[71][35] = 0;rain_draw[72][35] = 0;rain_draw[73][35] = 0;rain_draw[74][35] = 0;rain_draw[75][35] = 0;rain_draw[76][35] = 0;rain_draw[77][35] = 0;rain_draw[78][35] = 0;rain_draw[79][35] = 0;rain_draw[80][35] = 0;rain_draw[81][35] = 0;rain_draw[82][35] = 0;rain_draw[83][35] = 0;rain_draw[84][35] = 0;rain_draw[85][35] = 0;rain_draw[86][35] = 0;rain_draw[87][35] = 0;rain_draw[88][35] = 0;rain_draw[89][35] = 0;rain_draw[90][35] = 0;rain_draw[91][35] = 0;rain_draw[92][35] = 0;rain_draw[93][35] = 0;rain_draw[94][35] = 0;rain_draw[95][35] = 0;
        rain_draw[0][36] = 0;rain_draw[1][36] = 0;rain_draw[2][36] = 0;rain_draw[3][36] = 0;rain_draw[4][36] = 0;rain_draw[5][36] = 0;rain_draw[6][36] = 0;rain_draw[7][36] = 0;rain_draw[8][36] = 0;rain_draw[9][36] = 0;rain_draw[10][36] = 0;rain_draw[11][36] = 0;rain_draw[12][36] = 0;rain_draw[13][36] = 0;rain_draw[14][36] = 0;rain_draw[15][36] = 0;rain_draw[16][36] = 0;rain_draw[17][36] = 0;rain_draw[18][36] = 0;rain_draw[19][36] = 0;rain_draw[20][36] = 0;rain_draw[21][36] = 0;rain_draw[22][36] = 0;rain_draw[23][36] = 0;rain_draw[24][36] = 0;rain_draw[25][36] = 0;rain_draw[26][36] = 0;rain_draw[27][36] = 0;rain_draw[28][36] = 0;rain_draw[29][36] = 0;rain_draw[30][36] = 0;rain_draw[31][36] = 0;rain_draw[32][36] = 0;rain_draw[33][36] = 0;rain_draw[34][36] = 0;rain_draw[35][36] = 0;rain_draw[36][36] = 0;rain_draw[37][36] = 0;rain_draw[38][36] = 0;rain_draw[39][36] = 0;rain_draw[40][36] = 0;rain_draw[41][36] = 0;rain_draw[42][36] = 0;rain_draw[43][36] = 0;rain_draw[44][36] = 0;rain_draw[45][36] = 0;rain_draw[46][36] = 0;rain_draw[47][36] = 0;rain_draw[48][36] = 0;rain_draw[49][36] = 0;rain_draw[50][36] = 0;rain_draw[51][36] = 0;rain_draw[52][36] = 0;rain_draw[53][36] = 0;rain_draw[54][36] = 0;rain_draw[55][36] = 0;rain_draw[56][36] = 0;rain_draw[57][36] = 0;rain_draw[58][36] = 0;rain_draw[59][36] = 0;rain_draw[60][36] = 0;rain_draw[61][36] = 0;rain_draw[62][36] = 0;rain_draw[63][36] = 0;rain_draw[64][36] = 0;rain_draw[65][36] = 0;rain_draw[66][36] = 0;rain_draw[67][36] = 0;rain_draw[68][36] = 0;rain_draw[69][36] = 0;rain_draw[70][36] = 0;rain_draw[71][36] = 0;rain_draw[72][36] = 0;rain_draw[73][36] = 0;rain_draw[74][36] = 0;rain_draw[75][36] = 0;rain_draw[76][36] = 0;rain_draw[77][36] = 0;rain_draw[78][36] = 0;rain_draw[79][36] = 0;rain_draw[80][36] = 0;rain_draw[81][36] = 0;rain_draw[82][36] = 1;rain_draw[83][36] = 1;rain_draw[84][36] = 1;rain_draw[85][36] = 0;rain_draw[86][36] = 0;rain_draw[87][36] = 0;rain_draw[88][36] = 0;rain_draw[89][36] = 0;rain_draw[90][36] = 0;rain_draw[91][36] = 0;rain_draw[92][36] = 0;rain_draw[93][36] = 0;rain_draw[94][36] = 0;rain_draw[95][36] = 0;
        rain_draw[0][37] = 0;rain_draw[1][37] = 0;rain_draw[2][37] = 0;rain_draw[3][37] = 0;rain_draw[4][37] = 0;rain_draw[5][37] = 0;rain_draw[6][37] = 0;rain_draw[7][37] = 0;rain_draw[8][37] = 0;rain_draw[9][37] = 0;rain_draw[10][37] = 0;rain_draw[11][37] = 0;rain_draw[12][37] = 0;rain_draw[13][37] = 0;rain_draw[14][37] = 0;rain_draw[15][37] = 0;rain_draw[16][37] = 0;rain_draw[17][37] = 0;rain_draw[18][37] = 0;rain_draw[19][37] = 0;rain_draw[20][37] = 0;rain_draw[21][37] = 0;rain_draw[22][37] = 0;rain_draw[23][37] = 0;rain_draw[24][37] = 0;rain_draw[25][37] = 0;rain_draw[26][37] = 0;rain_draw[27][37] = 0;rain_draw[28][37] = 0;rain_draw[29][37] = 0;rain_draw[30][37] = 0;rain_draw[31][37] = 0;rain_draw[32][37] = 0;rain_draw[33][37] = 0;rain_draw[34][37] = 0;rain_draw[35][37] = 0;rain_draw[36][37] = 0;rain_draw[37][37] = 0;rain_draw[38][37] = 0;rain_draw[39][37] = 0;rain_draw[40][37] = 0;rain_draw[41][37] = 0;rain_draw[42][37] = 0;rain_draw[43][37] = 0;rain_draw[44][37] = 0;rain_draw[45][37] = 0;rain_draw[46][37] = 0;rain_draw[47][37] = 0;rain_draw[48][37] = 0;rain_draw[49][37] = 0;rain_draw[50][37] = 0;rain_draw[51][37] = 0;rain_draw[52][37] = 0;rain_draw[53][37] = 0;rain_draw[54][37] = 0;rain_draw[55][37] = 0;rain_draw[56][37] = 0;rain_draw[57][37] = 0;rain_draw[58][37] = 0;rain_draw[59][37] = 0;rain_draw[60][37] = 0;rain_draw[61][37] = 0;rain_draw[62][37] = 0;rain_draw[63][37] = 0;rain_draw[64][37] = 0;rain_draw[65][37] = 0;rain_draw[66][37] = 0;rain_draw[67][37] = 0;rain_draw[68][37] = 0;rain_draw[69][37] = 0;rain_draw[70][37] = 0;rain_draw[71][37] = 0;rain_draw[72][37] = 0;rain_draw[73][37] = 0;rain_draw[74][37] = 0;rain_draw[75][37] = 0;rain_draw[76][37] = 0;rain_draw[77][37] = 0;rain_draw[78][37] = 0;rain_draw[79][37] = 0;rain_draw[80][37] = 0;rain_draw[81][37] = 1;rain_draw[82][37] = 1;rain_draw[83][37] = 1;rain_draw[84][37] = 0;rain_draw[85][37] = 0;rain_draw[86][37] = 0;rain_draw[87][37] = 0;rain_draw[88][37] = 0;rain_draw[89][37] = 0;rain_draw[90][37] = 0;rain_draw[91][37] = 0;rain_draw[92][37] = 0;rain_draw[93][37] = 0;rain_draw[94][37] = 0;rain_draw[95][37] = 0;
        rain_draw[0][38] = 0;rain_draw[1][38] = 0;rain_draw[2][38] = 0;rain_draw[3][38] = 0;rain_draw[4][38] = 0;rain_draw[5][38] = 0;rain_draw[6][38] = 0;rain_draw[7][38] = 0;rain_draw[8][38] = 0;rain_draw[9][38] = 0;rain_draw[10][38] = 0;rain_draw[11][38] = 0;rain_draw[12][38] = 0;rain_draw[13][38] = 0;rain_draw[14][38] = 0;rain_draw[15][38] = 0;rain_draw[16][38] = 0;rain_draw[17][38] = 0;rain_draw[18][38] = 0;rain_draw[19][38] = 0;rain_draw[20][38] = 0;rain_draw[21][38] = 0;rain_draw[22][38] = 0;rain_draw[23][38] = 0;rain_draw[24][38] = 0;rain_draw[25][38] = 0;rain_draw[26][38] = 0;rain_draw[27][38] = 0;rain_draw[28][38] = 0;rain_draw[29][38] = 0;rain_draw[30][38] = 0;rain_draw[31][38] = 0;rain_draw[32][38] = 0;rain_draw[33][38] = 0;rain_draw[34][38] = 0;rain_draw[35][38] = 0;rain_draw[36][38] = 0;rain_draw[37][38] = 0;rain_draw[38][38] = 0;rain_draw[39][38] = 0;rain_draw[40][38] = 0;rain_draw[41][38] = 0;rain_draw[42][38] = 0;rain_draw[43][38] = 0;rain_draw[44][38] = 0;rain_draw[45][38] = 0;rain_draw[46][38] = 0;rain_draw[47][38] = 0;rain_draw[48][38] = 0;rain_draw[49][38] = 0;rain_draw[50][38] = 0;rain_draw[51][38] = 0;rain_draw[52][38] = 0;rain_draw[53][38] = 0;rain_draw[54][38] = 0;rain_draw[55][38] = 0;rain_draw[56][38] = 0;rain_draw[57][38] = 0;rain_draw[58][38] = 0;rain_draw[59][38] = 0;rain_draw[60][38] = 0;rain_draw[61][38] = 0;rain_draw[62][38] = 0;rain_draw[63][38] = 0;rain_draw[64][38] = 0;rain_draw[65][38] = 0;rain_draw[66][38] = 0;rain_draw[67][38] = 0;rain_draw[68][38] = 0;rain_draw[69][38] = 0;rain_draw[70][38] = 0;rain_draw[71][38] = 0;rain_draw[72][38] = 0;rain_draw[73][38] = 0;rain_draw[74][38] = 0;rain_draw[75][38] = 0;rain_draw[76][38] = 0;rain_draw[77][38] = 0;rain_draw[78][38] = 0;rain_draw[79][38] = 0;rain_draw[80][38] = 1;rain_draw[81][38] = 1;rain_draw[82][38] = 1;rain_draw[83][38] = 0;rain_draw[84][38] = 0;rain_draw[85][38] = 0;rain_draw[86][38] = 0;rain_draw[87][38] = 0;rain_draw[88][38] = 0;rain_draw[89][38] = 0;rain_draw[90][38] = 0;rain_draw[91][38] = 0;rain_draw[92][38] = 0;rain_draw[93][38] = 0;rain_draw[94][38] = 0;rain_draw[95][38] = 0;
        rain_draw[0][39] = 0;rain_draw[1][39] = 0;rain_draw[2][39] = 0;rain_draw[3][39] = 0;rain_draw[4][39] = 0;rain_draw[5][39] = 0;rain_draw[6][39] = 0;rain_draw[7][39] = 0;rain_draw[8][39] = 0;rain_draw[9][39] = 0;rain_draw[10][39] = 0;rain_draw[11][39] = 0;rain_draw[12][39] = 0;rain_draw[13][39] = 0;rain_draw[14][39] = 0;rain_draw[15][39] = 0;rain_draw[16][39] = 0;rain_draw[17][39] = 0;rain_draw[18][39] = 0;rain_draw[19][39] = 0;rain_draw[20][39] = 0;rain_draw[21][39] = 0;rain_draw[22][39] = 0;rain_draw[23][39] = 0;rain_draw[24][39] = 0;rain_draw[25][39] = 0;rain_draw[26][39] = 0;rain_draw[27][39] = 0;rain_draw[28][39] = 0;rain_draw[29][39] = 0;rain_draw[30][39] = 0;rain_draw[31][39] = 0;rain_draw[32][39] = 0;rain_draw[33][39] = 0;rain_draw[34][39] = 0;rain_draw[35][39] = 0;rain_draw[36][39] = 0;rain_draw[37][39] = 0;rain_draw[38][39] = 0;rain_draw[39][39] = 0;rain_draw[40][39] = 0;rain_draw[41][39] = 0;rain_draw[42][39] = 0;rain_draw[43][39] = 0;rain_draw[44][39] = 0;rain_draw[45][39] = 0;rain_draw[46][39] = 0;rain_draw[47][39] = 0;rain_draw[48][39] = 0;rain_draw[49][39] = 0;rain_draw[50][39] = 0;rain_draw[51][39] = 0;rain_draw[52][39] = 0;rain_draw[53][39] = 0;rain_draw[54][39] = 0;rain_draw[55][39] = 0;rain_draw[56][39] = 0;rain_draw[57][39] = 0;rain_draw[58][39] = 0;rain_draw[59][39] = 0;rain_draw[60][39] = 0;rain_draw[61][39] = 0;rain_draw[62][39] = 0;rain_draw[63][39] = 0;rain_draw[64][39] = 0;rain_draw[65][39] = 0;rain_draw[66][39] = 0;rain_draw[67][39] = 0;rain_draw[68][39] = 0;rain_draw[69][39] = 0;rain_draw[70][39] = 0;rain_draw[71][39] = 0;rain_draw[72][39] = 0;rain_draw[73][39] = 0;rain_draw[74][39] = 0;rain_draw[75][39] = 0;rain_draw[76][39] = 0;rain_draw[77][39] = 0;rain_draw[78][39] = 0;rain_draw[79][39] = 1;rain_draw[80][39] = 1;rain_draw[81][39] = 1;rain_draw[82][39] = 0;rain_draw[83][39] = 0;rain_draw[84][39] = 0;rain_draw[85][39] = 0;rain_draw[86][39] = 0;rain_draw[87][39] = 0;rain_draw[88][39] = 0;rain_draw[89][39] = 0;rain_draw[90][39] = 0;rain_draw[91][39] = 0;rain_draw[92][39] = 0;rain_draw[93][39] = 0;rain_draw[94][39] = 0;rain_draw[95][39] = 0;
        rain_draw[0][40] = 0;rain_draw[1][40] = 0;rain_draw[2][40] = 0;rain_draw[3][40] = 0;rain_draw[4][40] = 0;rain_draw[5][40] = 0;rain_draw[6][40] = 0;rain_draw[7][40] = 0;rain_draw[8][40] = 0;rain_draw[9][40] = 0;rain_draw[10][40] = 0;rain_draw[11][40] = 0;rain_draw[12][40] = 0;rain_draw[13][40] = 0;rain_draw[14][40] = 0;rain_draw[15][40] = 0;rain_draw[16][40] = 0;rain_draw[17][40] = 0;rain_draw[18][40] = 0;rain_draw[19][40] = 0;rain_draw[20][40] = 0;rain_draw[21][40] = 0;rain_draw[22][40] = 0;rain_draw[23][40] = 0;rain_draw[24][40] = 0;rain_draw[25][40] = 0;rain_draw[26][40] = 0;rain_draw[27][40] = 0;rain_draw[28][40] = 0;rain_draw[29][40] = 0;rain_draw[30][40] = 0;rain_draw[31][40] = 0;rain_draw[32][40] = 0;rain_draw[33][40] = 0;rain_draw[34][40] = 0;rain_draw[35][40] = 0;rain_draw[36][40] = 0;rain_draw[37][40] = 0;rain_draw[38][40] = 0;rain_draw[39][40] = 0;rain_draw[40][40] = 0;rain_draw[41][40] = 0;rain_draw[42][40] = 0;rain_draw[43][40] = 0;rain_draw[44][40] = 0;rain_draw[45][40] = 0;rain_draw[46][40] = 0;rain_draw[47][40] = 0;rain_draw[48][40] = 0;rain_draw[49][40] = 0;rain_draw[50][40] = 0;rain_draw[51][40] = 0;rain_draw[52][40] = 0;rain_draw[53][40] = 0;rain_draw[54][40] = 0;rain_draw[55][40] = 0;rain_draw[56][40] = 0;rain_draw[57][40] = 0;rain_draw[58][40] = 0;rain_draw[59][40] = 0;rain_draw[60][40] = 0;rain_draw[61][40] = 0;rain_draw[62][40] = 0;rain_draw[63][40] = 0;rain_draw[64][40] = 0;rain_draw[65][40] = 0;rain_draw[66][40] = 0;rain_draw[67][40] = 0;rain_draw[68][40] = 0;rain_draw[69][40] = 0;rain_draw[70][40] = 0;rain_draw[71][40] = 0;rain_draw[72][40] = 0;rain_draw[73][40] = 0;rain_draw[74][40] = 0;rain_draw[75][40] = 0;rain_draw[76][40] = 0;rain_draw[77][40] = 0;rain_draw[78][40] = 1;rain_draw[79][40] = 1;rain_draw[80][40] = 1;rain_draw[81][40] = 0;rain_draw[82][40] = 0;rain_draw[83][40] = 0;rain_draw[84][40] = 0;rain_draw[85][40] = 0;rain_draw[86][40] = 0;rain_draw[87][40] = 0;rain_draw[88][40] = 0;rain_draw[89][40] = 0;rain_draw[90][40] = 0;rain_draw[91][40] = 0;rain_draw[92][40] = 0;rain_draw[93][40] = 0;rain_draw[94][40] = 0;rain_draw[95][40] = 0;
        rain_draw[0][41] = 0;rain_draw[1][41] = 0;rain_draw[2][41] = 0;rain_draw[3][41] = 0;rain_draw[4][41] = 0;rain_draw[5][41] = 0;rain_draw[6][41] = 0;rain_draw[7][41] = 0;rain_draw[8][41] = 0;rain_draw[9][41] = 0;rain_draw[10][41] = 0;rain_draw[11][41] = 0;rain_draw[12][41] = 0;rain_draw[13][41] = 0;rain_draw[14][41] = 0;rain_draw[15][41] = 0;rain_draw[16][41] = 0;rain_draw[17][41] = 0;rain_draw[18][41] = 0;rain_draw[19][41] = 0;rain_draw[20][41] = 0;rain_draw[21][41] = 0;rain_draw[22][41] = 0;rain_draw[23][41] = 0;rain_draw[24][41] = 0;rain_draw[25][41] = 0;rain_draw[26][41] = 0;rain_draw[27][41] = 0;rain_draw[28][41] = 0;rain_draw[29][41] = 1;rain_draw[30][41] = 1;rain_draw[31][41] = 1;rain_draw[32][41] = 0;rain_draw[33][41] = 0;rain_draw[34][41] = 0;rain_draw[35][41] = 0;rain_draw[36][41] = 0;rain_draw[37][41] = 0;rain_draw[38][41] = 0;rain_draw[39][41] = 0;rain_draw[40][41] = 0;rain_draw[41][41] = 0;rain_draw[42][41] = 0;rain_draw[43][41] = 0;rain_draw[44][41] = 0;rain_draw[45][41] = 0;rain_draw[46][41] = 0;rain_draw[47][41] = 0;rain_draw[48][41] = 0;rain_draw[49][41] = 0;rain_draw[50][41] = 0;rain_draw[51][41] = 0;rain_draw[52][41] = 0;rain_draw[53][41] = 0;rain_draw[54][41] = 0;rain_draw[55][41] = 0;rain_draw[56][41] = 0;rain_draw[57][41] = 0;rain_draw[58][41] = 0;rain_draw[59][41] = 0;rain_draw[60][41] = 0;rain_draw[61][41] = 0;rain_draw[62][41] = 0;rain_draw[63][41] = 0;rain_draw[64][41] = 0;rain_draw[65][41] = 0;rain_draw[66][41] = 0;rain_draw[67][41] = 0;rain_draw[68][41] = 0;rain_draw[69][41] = 0;rain_draw[70][41] = 0;rain_draw[71][41] = 0;rain_draw[72][41] = 0;rain_draw[73][41] = 0;rain_draw[74][41] = 0;rain_draw[75][41] = 0;rain_draw[76][41] = 0;rain_draw[77][41] = 1;rain_draw[78][41] = 1;rain_draw[79][41] = 1;rain_draw[80][41] = 0;rain_draw[81][41] = 0;rain_draw[82][41] = 0;rain_draw[83][41] = 0;rain_draw[84][41] = 0;rain_draw[85][41] = 0;rain_draw[86][41] = 0;rain_draw[87][41] = 0;rain_draw[88][41] = 0;rain_draw[89][41] = 0;rain_draw[90][41] = 0;rain_draw[91][41] = 0;rain_draw[92][41] = 0;rain_draw[93][41] = 0;rain_draw[94][41] = 0;rain_draw[95][41] = 0;
        rain_draw[0][42] = 0;rain_draw[1][42] = 0;rain_draw[2][42] = 0;rain_draw[3][42] = 0;rain_draw[4][42] = 0;rain_draw[5][42] = 0;rain_draw[6][42] = 0;rain_draw[7][42] = 0;rain_draw[8][42] = 0;rain_draw[9][42] = 0;rain_draw[10][42] = 0;rain_draw[11][42] = 0;rain_draw[12][42] = 0;rain_draw[13][42] = 0;rain_draw[14][42] = 0;rain_draw[15][42] = 0;rain_draw[16][42] = 0;rain_draw[17][42] = 0;rain_draw[18][42] = 0;rain_draw[19][42] = 0;rain_draw[20][42] = 0;rain_draw[21][42] = 0;rain_draw[22][42] = 0;rain_draw[23][42] = 0;rain_draw[24][42] = 0;rain_draw[25][42] = 0;rain_draw[26][42] = 0;rain_draw[27][42] = 0;rain_draw[28][42] = 1;rain_draw[29][42] = 1;rain_draw[30][42] = 1;rain_draw[31][42] = 0;rain_draw[32][42] = 0;rain_draw[33][42] = 0;rain_draw[34][42] = 0;rain_draw[35][42] = 0;rain_draw[36][42] = 0;rain_draw[37][42] = 0;rain_draw[38][42] = 0;rain_draw[39][42] = 0;rain_draw[40][42] = 0;rain_draw[41][42] = 0;rain_draw[42][42] = 0;rain_draw[43][42] = 0;rain_draw[44][42] = 0;rain_draw[45][42] = 0;rain_draw[46][42] = 0;rain_draw[47][42] = 0;rain_draw[48][42] = 0;rain_draw[49][42] = 0;rain_draw[50][42] = 0;rain_draw[51][42] = 0;rain_draw[52][42] = 0;rain_draw[53][42] = 0;rain_draw[54][42] = 0;rain_draw[55][42] = 0;rain_draw[56][42] = 0;rain_draw[57][42] = 0;rain_draw[58][42] = 0;rain_draw[59][42] = 0;rain_draw[60][42] = 0;rain_draw[61][42] = 0;rain_draw[62][42] = 0;rain_draw[63][42] = 0;rain_draw[64][42] = 0;rain_draw[65][42] = 0;rain_draw[66][42] = 0;rain_draw[67][42] = 0;rain_draw[68][42] = 0;rain_draw[69][42] = 0;rain_draw[70][42] = 0;rain_draw[71][42] = 0;rain_draw[72][42] = 0;rain_draw[73][42] = 0;rain_draw[74][42] = 0;rain_draw[75][42] = 0;rain_draw[76][42] = 1;rain_draw[77][42] = 1;rain_draw[78][42] = 1;rain_draw[79][42] = 0;rain_draw[80][42] = 0;rain_draw[81][42] = 0;rain_draw[82][42] = 0;rain_draw[83][42] = 0;rain_draw[84][42] = 0;rain_draw[85][42] = 0;rain_draw[86][42] = 0;rain_draw[87][42] = 0;rain_draw[88][42] = 0;rain_draw[89][42] = 0;rain_draw[90][42] = 0;rain_draw[91][42] = 0;rain_draw[92][42] = 0;rain_draw[93][42] = 0;rain_draw[94][42] = 0;rain_draw[95][42] = 0;
        rain_draw[0][43] = 0;rain_draw[1][43] = 0;rain_draw[2][43] = 0;rain_draw[3][43] = 0;rain_draw[4][43] = 0;rain_draw[5][43] = 0;rain_draw[6][43] = 0;rain_draw[7][43] = 0;rain_draw[8][43] = 0;rain_draw[9][43] = 0;rain_draw[10][43] = 0;rain_draw[11][43] = 0;rain_draw[12][43] = 0;rain_draw[13][43] = 0;rain_draw[14][43] = 0;rain_draw[15][43] = 0;rain_draw[16][43] = 0;rain_draw[17][43] = 0;rain_draw[18][43] = 0;rain_draw[19][43] = 0;rain_draw[20][43] = 0;rain_draw[21][43] = 0;rain_draw[22][43] = 0;rain_draw[23][43] = 0;rain_draw[24][43] = 0;rain_draw[25][43] = 0;rain_draw[26][43] = 0;rain_draw[27][43] = 1;rain_draw[28][43] = 1;rain_draw[29][43] = 1;rain_draw[30][43] = 0;rain_draw[31][43] = 0;rain_draw[32][43] = 0;rain_draw[33][43] = 0;rain_draw[34][43] = 0;rain_draw[35][43] = 0;rain_draw[36][43] = 0;rain_draw[37][43] = 0;rain_draw[38][43] = 0;rain_draw[39][43] = 0;rain_draw[40][43] = 0;rain_draw[41][43] = 0;rain_draw[42][43] = 0;rain_draw[43][43] = 0;rain_draw[44][43] = 0;rain_draw[45][43] = 0;rain_draw[46][43] = 0;rain_draw[47][43] = 0;rain_draw[48][43] = 0;rain_draw[49][43] = 0;rain_draw[50][43] = 0;rain_draw[51][43] = 0;rain_draw[52][43] = 0;rain_draw[53][43] = 0;rain_draw[54][43] = 0;rain_draw[55][43] = 0;rain_draw[56][43] = 0;rain_draw[57][43] = 0;rain_draw[58][43] = 0;rain_draw[59][43] = 0;rain_draw[60][43] = 0;rain_draw[61][43] = 0;rain_draw[62][43] = 0;rain_draw[63][43] = 0;rain_draw[64][43] = 0;rain_draw[65][43] = 0;rain_draw[66][43] = 0;rain_draw[67][43] = 0;rain_draw[68][43] = 0;rain_draw[69][43] = 0;rain_draw[70][43] = 0;rain_draw[71][43] = 0;rain_draw[72][43] = 0;rain_draw[73][43] = 0;rain_draw[74][43] = 0;rain_draw[75][43] = 0;rain_draw[76][43] = 0;rain_draw[77][43] = 0;rain_draw[78][43] = 0;rain_draw[79][43] = 0;rain_draw[80][43] = 0;rain_draw[81][43] = 0;rain_draw[82][43] = 0;rain_draw[83][43] = 0;rain_draw[84][43] = 0;rain_draw[85][43] = 0;rain_draw[86][43] = 0;rain_draw[87][43] = 0;rain_draw[88][43] = 0;rain_draw[89][43] = 0;rain_draw[90][43] = 0;rain_draw[91][43] = 0;rain_draw[92][43] = 0;rain_draw[93][43] = 0;rain_draw[94][43] = 0;rain_draw[95][43] = 0;
        rain_draw[0][44] = 0;rain_draw[1][44] = 0;rain_draw[2][44] = 0;rain_draw[3][44] = 0;rain_draw[4][44] = 0;rain_draw[5][44] = 0;rain_draw[6][44] = 0;rain_draw[7][44] = 0;rain_draw[8][44] = 0;rain_draw[9][44] = 1;rain_draw[10][44] = 1;rain_draw[11][44] = 1;rain_draw[12][44] = 0;rain_draw[13][44] = 0;rain_draw[14][44] = 0;rain_draw[15][44] = 0;rain_draw[16][44] = 0;rain_draw[17][44] = 0;rain_draw[18][44] = 0;rain_draw[19][44] = 0;rain_draw[20][44] = 0;rain_draw[21][44] = 0;rain_draw[22][44] = 0;rain_draw[23][44] = 0;rain_draw[24][44] = 0;rain_draw[25][44] = 0;rain_draw[26][44] = 1;rain_draw[27][44] = 1;rain_draw[28][44] = 1;rain_draw[29][44] = 0;rain_draw[30][44] = 0;rain_draw[31][44] = 0;rain_draw[32][44] = 0;rain_draw[33][44] = 0;rain_draw[34][44] = 0;rain_draw[35][44] = 0;rain_draw[36][44] = 0;rain_draw[37][44] = 0;rain_draw[38][44] = 0;rain_draw[39][44] = 0;rain_draw[40][44] = 0;rain_draw[41][44] = 0;rain_draw[42][44] = 0;rain_draw[43][44] = 0;rain_draw[44][44] = 0;rain_draw[45][44] = 0;rain_draw[46][44] = 0;rain_draw[47][44] = 0;rain_draw[48][44] = 0;rain_draw[49][44] = 0;rain_draw[50][44] = 0;rain_draw[51][44] = 0;rain_draw[52][44] = 0;rain_draw[53][44] = 0;rain_draw[54][44] = 0;rain_draw[55][44] = 0;rain_draw[56][44] = 0;rain_draw[57][44] = 0;rain_draw[58][44] = 0;rain_draw[59][44] = 0;rain_draw[60][44] = 0;rain_draw[61][44] = 0;rain_draw[62][44] = 0;rain_draw[63][44] = 0;rain_draw[64][44] = 0;rain_draw[65][44] = 0;rain_draw[66][44] = 0;rain_draw[67][44] = 0;rain_draw[68][44] = 0;rain_draw[69][44] = 0;rain_draw[70][44] = 0;rain_draw[71][44] = 0;rain_draw[72][44] = 0;rain_draw[73][44] = 0;rain_draw[74][44] = 0;rain_draw[75][44] = 0;rain_draw[76][44] = 0;rain_draw[77][44] = 0;rain_draw[78][44] = 0;rain_draw[79][44] = 0;rain_draw[80][44] = 0;rain_draw[81][44] = 0;rain_draw[82][44] = 0;rain_draw[83][44] = 0;rain_draw[84][44] = 0;rain_draw[85][44] = 0;rain_draw[86][44] = 0;rain_draw[87][44] = 0;rain_draw[88][44] = 0;rain_draw[89][44] = 0;rain_draw[90][44] = 0;rain_draw[91][44] = 0;rain_draw[92][44] = 0;rain_draw[93][44] = 0;rain_draw[94][44] = 0;rain_draw[95][44] = 0;
        rain_draw[0][45] = 0;rain_draw[1][45] = 0;rain_draw[2][45] = 0;rain_draw[3][45] = 0;rain_draw[4][45] = 0;rain_draw[5][45] = 0;rain_draw[6][45] = 0;rain_draw[7][45] = 0;rain_draw[8][45] = 1;rain_draw[9][45] = 1;rain_draw[10][45] = 1;rain_draw[11][45] = 0;rain_draw[12][45] = 0;rain_draw[13][45] = 0;rain_draw[14][45] = 0;rain_draw[15][45] = 0;rain_draw[16][45] = 0;rain_draw[17][45] = 0;rain_draw[18][45] = 0;rain_draw[19][45] = 0;rain_draw[20][45] = 0;rain_draw[21][45] = 0;rain_draw[22][45] = 0;rain_draw[23][45] = 0;rain_draw[24][45] = 0;rain_draw[25][45] = 1;rain_draw[26][45] = 1;rain_draw[27][45] = 1;rain_draw[28][45] = 0;rain_draw[29][45] = 0;rain_draw[30][45] = 0;rain_draw[31][45] = 0;rain_draw[32][45] = 0;rain_draw[33][45] = 0;rain_draw[34][45] = 0;rain_draw[35][45] = 0;rain_draw[36][45] = 0;rain_draw[37][45] = 0;rain_draw[38][45] = 0;rain_draw[39][45] = 0;rain_draw[40][45] = 0;rain_draw[41][45] = 0;rain_draw[42][45] = 0;rain_draw[43][45] = 0;rain_draw[44][45] = 0;rain_draw[45][45] = 0;rain_draw[46][45] = 0;rain_draw[47][45] = 0;rain_draw[48][45] = 0;rain_draw[49][45] = 0;rain_draw[50][45] = 0;rain_draw[51][45] = 0;rain_draw[52][45] = 0;rain_draw[53][45] = 0;rain_draw[54][45] = 0;rain_draw[55][45] = 0;rain_draw[56][45] = 0;rain_draw[57][45] = 0;rain_draw[58][45] = 0;rain_draw[59][45] = 0;rain_draw[60][45] = 0;rain_draw[61][45] = 0;rain_draw[62][45] = 0;rain_draw[63][45] = 0;rain_draw[64][45] = 0;rain_draw[65][45] = 0;rain_draw[66][45] = 0;rain_draw[67][45] = 0;rain_draw[68][45] = 0;rain_draw[69][45] = 0;rain_draw[70][45] = 0;rain_draw[71][45] = 0;rain_draw[72][45] = 0;rain_draw[73][45] = 0;rain_draw[74][45] = 0;rain_draw[75][45] = 0;rain_draw[76][45] = 0;rain_draw[77][45] = 0;rain_draw[78][45] = 0;rain_draw[79][45] = 0;rain_draw[80][45] = 0;rain_draw[81][45] = 0;rain_draw[82][45] = 0;rain_draw[83][45] = 0;rain_draw[84][45] = 0;rain_draw[85][45] = 0;rain_draw[86][45] = 0;rain_draw[87][45] = 0;rain_draw[88][45] = 0;rain_draw[89][45] = 0;rain_draw[90][45] = 0;rain_draw[91][45] = 0;rain_draw[92][45] = 0;rain_draw[93][45] = 0;rain_draw[94][45] = 0;rain_draw[95][45] = 0;
        rain_draw[0][46] = 0;rain_draw[1][46] = 0;rain_draw[2][46] = 0;rain_draw[3][46] = 0;rain_draw[4][46] = 0;rain_draw[5][46] = 0;rain_draw[6][46] = 0;rain_draw[7][46] = 1;rain_draw[8][46] = 1;rain_draw[9][46] = 1;rain_draw[10][46] = 0;rain_draw[11][46] = 0;rain_draw[12][46] = 0;rain_draw[13][46] = 0;rain_draw[14][46] = 0;rain_draw[15][46] = 0;rain_draw[16][46] = 0;rain_draw[17][46] = 0;rain_draw[18][46] = 0;rain_draw[19][46] = 0;rain_draw[20][46] = 0;rain_draw[21][46] = 0;rain_draw[22][46] = 0;rain_draw[23][46] = 0;rain_draw[24][46] = 1;rain_draw[25][46] = 1;rain_draw[26][46] = 1;rain_draw[27][46] = 0;rain_draw[28][46] = 0;rain_draw[29][46] = 0;rain_draw[30][46] = 0;rain_draw[31][46] = 0;rain_draw[32][46] = 0;rain_draw[33][46] = 0;rain_draw[34][46] = 0;rain_draw[35][46] = 0;rain_draw[36][46] = 0;rain_draw[37][46] = 0;rain_draw[38][46] = 0;rain_draw[39][46] = 0;rain_draw[40][46] = 0;rain_draw[41][46] = 1;rain_draw[42][46] = 1;rain_draw[43][46] = 1;rain_draw[44][46] = 0;rain_draw[45][46] = 0;rain_draw[46][46] = 0;rain_draw[47][46] = 0;rain_draw[48][46] = 0;rain_draw[49][46] = 0;rain_draw[50][46] = 0;rain_draw[51][46] = 0;rain_draw[52][46] = 0;rain_draw[53][46] = 0;rain_draw[54][46] = 0;rain_draw[55][46] = 0;rain_draw[56][46] = 0;rain_draw[57][46] = 0;rain_draw[58][46] = 0;rain_draw[59][46] = 0;rain_draw[60][46] = 0;rain_draw[61][46] = 0;rain_draw[62][46] = 0;rain_draw[63][46] = 0;rain_draw[64][46] = 0;rain_draw[65][46] = 0;rain_draw[66][46] = 0;rain_draw[67][46] = 0;rain_draw[68][46] = 0;rain_draw[69][46] = 0;rain_draw[70][46] = 0;rain_draw[71][46] = 0;rain_draw[72][46] = 0;rain_draw[73][46] = 0;rain_draw[74][46] = 0;rain_draw[75][46] = 0;rain_draw[76][46] = 0;rain_draw[77][46] = 0;rain_draw[78][46] = 0;rain_draw[79][46] = 0;rain_draw[80][46] = 0;rain_draw[81][46] = 0;rain_draw[82][46] = 0;rain_draw[83][46] = 0;rain_draw[84][46] = 0;rain_draw[85][46] = 0;rain_draw[86][46] = 0;rain_draw[87][46] = 0;rain_draw[88][46] = 0;rain_draw[89][46] = 0;rain_draw[90][46] = 0;rain_draw[91][46] = 0;rain_draw[92][46] = 0;rain_draw[93][46] = 0;rain_draw[94][46] = 0;rain_draw[95][46] = 0;
        rain_draw[0][47] = 0;rain_draw[1][47] = 0;rain_draw[2][47] = 0;rain_draw[3][47] = 0;rain_draw[4][47] = 0;rain_draw[5][47] = 0;rain_draw[6][47] = 1;rain_draw[7][47] = 1;rain_draw[8][47] = 1;rain_draw[9][47] = 0;rain_draw[10][47] = 0;rain_draw[11][47] = 0;rain_draw[12][47] = 0;rain_draw[13][47] = 0;rain_draw[14][47] = 0;rain_draw[15][47] = 0;rain_draw[16][47] = 0;rain_draw[17][47] = 0;rain_draw[18][47] = 0;rain_draw[19][47] = 0;rain_draw[20][47] = 0;rain_draw[21][47] = 0;rain_draw[22][47] = 0;rain_draw[23][47] = 1;rain_draw[24][47] = 1;rain_draw[25][47] = 1;rain_draw[26][47] = 0;rain_draw[27][47] = 0;rain_draw[28][47] = 0;rain_draw[29][47] = 0;rain_draw[30][47] = 0;rain_draw[31][47] = 0;rain_draw[32][47] = 0;rain_draw[33][47] = 0;rain_draw[34][47] = 0;rain_draw[35][47] = 0;rain_draw[36][47] = 0;rain_draw[37][47] = 0;rain_draw[38][47] = 0;rain_draw[39][47] = 0;rain_draw[40][47] = 1;rain_draw[41][47] = 1;rain_draw[42][47] = 1;rain_draw[43][47] = 0;rain_draw[44][47] = 0;rain_draw[45][47] = 0;rain_draw[46][47] = 0;rain_draw[47][47] = 0;rain_draw[48][47] = 0;rain_draw[49][47] = 0;rain_draw[50][47] = 0;rain_draw[51][47] = 0;rain_draw[52][47] = 0;rain_draw[53][47] = 0;rain_draw[54][47] = 0;rain_draw[55][47] = 0;rain_draw[56][47] = 0;rain_draw[57][47] = 0;rain_draw[58][47] = 0;rain_draw[59][47] = 0;rain_draw[60][47] = 0;rain_draw[61][47] = 0;rain_draw[62][47] = 0;rain_draw[63][47] = 0;rain_draw[64][47] = 0;rain_draw[65][47] = 0;rain_draw[66][47] = 0;rain_draw[67][47] = 0;rain_draw[68][47] = 0;rain_draw[69][47] = 0;rain_draw[70][47] = 0;rain_draw[71][47] = 0;rain_draw[72][47] = 0;rain_draw[73][47] = 0;rain_draw[74][47] = 0;rain_draw[75][47] = 0;rain_draw[76][47] = 0;rain_draw[77][47] = 0;rain_draw[78][47] = 0;rain_draw[79][47] = 0;rain_draw[80][47] = 0;rain_draw[81][47] = 0;rain_draw[82][47] = 0;rain_draw[83][47] = 0;rain_draw[84][47] = 0;rain_draw[85][47] = 0;rain_draw[86][47] = 0;rain_draw[87][47] = 0;rain_draw[88][47] = 0;rain_draw[89][47] = 0;rain_draw[90][47] = 0;rain_draw[91][47] = 0;rain_draw[92][47] = 0;rain_draw[93][47] = 0;rain_draw[94][47] = 0;rain_draw[95][47] = 0;
        rain_draw[0][48] = 0;rain_draw[1][48] = 0;rain_draw[2][48] = 0;rain_draw[3][48] = 0;rain_draw[4][48] = 0;rain_draw[5][48] = 1;rain_draw[6][48] = 1;rain_draw[7][48] = 1;rain_draw[8][48] = 0;rain_draw[9][48] = 0;rain_draw[10][48] = 0;rain_draw[11][48] = 0;rain_draw[12][48] = 0;rain_draw[13][48] = 0;rain_draw[14][48] = 0;rain_draw[15][48] = 0;rain_draw[16][48] = 0;rain_draw[17][48] = 0;rain_draw[18][48] = 0;rain_draw[19][48] = 0;rain_draw[20][48] = 0;rain_draw[21][48] = 0;rain_draw[22][48] = 0;rain_draw[23][48] = 0;rain_draw[24][48] = 0;rain_draw[25][48] = 0;rain_draw[26][48] = 0;rain_draw[27][48] = 0;rain_draw[28][48] = 0;rain_draw[29][48] = 0;rain_draw[30][48] = 0;rain_draw[31][48] = 0;rain_draw[32][48] = 0;rain_draw[33][48] = 0;rain_draw[34][48] = 0;rain_draw[35][48] = 0;rain_draw[36][48] = 0;rain_draw[37][48] = 0;rain_draw[38][48] = 0;rain_draw[39][48] = 1;rain_draw[40][48] = 1;rain_draw[41][48] = 1;rain_draw[42][48] = 0;rain_draw[43][48] = 0;rain_draw[44][48] = 0;rain_draw[45][48] = 0;rain_draw[46][48] = 0;rain_draw[47][48] = 0;rain_draw[48][48] = 0;rain_draw[49][48] = 0;rain_draw[50][48] = 0;rain_draw[51][48] = 0;rain_draw[52][48] = 0;rain_draw[53][48] = 0;rain_draw[54][48] = 0;rain_draw[55][48] = 0;rain_draw[56][48] = 0;rain_draw[57][48] = 0;rain_draw[58][48] = 0;rain_draw[59][48] = 0;rain_draw[60][48] = 0;rain_draw[61][48] = 0;rain_draw[62][48] = 0;rain_draw[63][48] = 0;rain_draw[64][48] = 0;rain_draw[65][48] = 0;rain_draw[66][48] = 0;rain_draw[67][48] = 0;rain_draw[68][48] = 0;rain_draw[69][48] = 0;rain_draw[70][48] = 0;rain_draw[71][48] = 0;rain_draw[72][48] = 0;rain_draw[73][48] = 0;rain_draw[74][48] = 0;rain_draw[75][48] = 0;rain_draw[76][48] = 0;rain_draw[77][48] = 0;rain_draw[78][48] = 0;rain_draw[79][48] = 0;rain_draw[80][48] = 0;rain_draw[81][48] = 0;rain_draw[82][48] = 0;rain_draw[83][48] = 0;rain_draw[84][48] = 0;rain_draw[85][48] = 0;rain_draw[86][48] = 0;rain_draw[87][48] = 0;rain_draw[88][48] = 0;rain_draw[89][48] = 0;rain_draw[90][48] = 0;rain_draw[91][48] = 0;rain_draw[92][48] = 0;rain_draw[93][48] = 0;rain_draw[94][48] = 0;rain_draw[95][48] = 0;
        rain_draw[0][49] = 0;rain_draw[1][49] = 0;rain_draw[2][49] = 0;rain_draw[3][49] = 0;rain_draw[4][49] = 1;rain_draw[5][49] = 1;rain_draw[6][49] = 1;rain_draw[7][49] = 0;rain_draw[8][49] = 0;rain_draw[9][49] = 0;rain_draw[10][49] = 0;rain_draw[11][49] = 0;rain_draw[12][49] = 0;rain_draw[13][49] = 0;rain_draw[14][49] = 0;rain_draw[15][49] = 0;rain_draw[16][49] = 0;rain_draw[17][49] = 0;rain_draw[18][49] = 0;rain_draw[19][49] = 0;rain_draw[20][49] = 0;rain_draw[21][49] = 0;rain_draw[22][49] = 0;rain_draw[23][49] = 0;rain_draw[24][49] = 0;rain_draw[25][49] = 0;rain_draw[26][49] = 0;rain_draw[27][49] = 0;rain_draw[28][49] = 0;rain_draw[29][49] = 0;rain_draw[30][49] = 0;rain_draw[31][49] = 0;rain_draw[32][49] = 0;rain_draw[33][49] = 0;rain_draw[34][49] = 0;rain_draw[35][49] = 0;rain_draw[36][49] = 0;rain_draw[37][49] = 0;rain_draw[38][49] = 1;rain_draw[39][49] = 1;rain_draw[40][49] = 1;rain_draw[41][49] = 0;rain_draw[42][49] = 0;rain_draw[43][49] = 0;rain_draw[44][49] = 0;rain_draw[45][49] = 0;rain_draw[46][49] = 0;rain_draw[47][49] = 0;rain_draw[48][49] = 0;rain_draw[49][49] = 0;rain_draw[50][49] = 0;rain_draw[51][49] = 0;rain_draw[52][49] = 0;rain_draw[53][49] = 0;rain_draw[54][49] = 0;rain_draw[55][49] = 0;rain_draw[56][49] = 0;rain_draw[57][49] = 0;rain_draw[58][49] = 0;rain_draw[59][49] = 0;rain_draw[60][49] = 0;rain_draw[61][49] = 0;rain_draw[62][49] = 0;rain_draw[63][49] = 0;rain_draw[64][49] = 0;rain_draw[65][49] = 0;rain_draw[66][49] = 0;rain_draw[67][49] = 0;rain_draw[68][49] = 0;rain_draw[69][49] = 0;rain_draw[70][49] = 0;rain_draw[71][49] = 0;rain_draw[72][49] = 0;rain_draw[73][49] = 0;rain_draw[74][49] = 0;rain_draw[75][49] = 0;rain_draw[76][49] = 0;rain_draw[77][49] = 0;rain_draw[78][49] = 0;rain_draw[79][49] = 0;rain_draw[80][49] = 0;rain_draw[81][49] = 0;rain_draw[82][49] = 0;rain_draw[83][49] = 0;rain_draw[84][49] = 0;rain_draw[85][49] = 0;rain_draw[86][49] = 0;rain_draw[87][49] = 0;rain_draw[88][49] = 0;rain_draw[89][49] = 0;rain_draw[90][49] = 0;rain_draw[91][49] = 0;rain_draw[92][49] = 0;rain_draw[93][49] = 0;rain_draw[94][49] = 0;rain_draw[95][49] = 0;
        rain_draw[0][50] = 0;rain_draw[1][50] = 0;rain_draw[2][50] = 0;rain_draw[3][50] = 1;rain_draw[4][50] = 1;rain_draw[5][50] = 1;rain_draw[6][50] = 0;rain_draw[7][50] = 0;rain_draw[8][50] = 0;rain_draw[9][50] = 0;rain_draw[10][50] = 0;rain_draw[11][50] = 0;rain_draw[12][50] = 0;rain_draw[13][50] = 0;rain_draw[14][50] = 0;rain_draw[15][50] = 0;rain_draw[16][50] = 0;rain_draw[17][50] = 0;rain_draw[18][50] = 0;rain_draw[19][50] = 0;rain_draw[20][50] = 0;rain_draw[21][50] = 0;rain_draw[22][50] = 0;rain_draw[23][50] = 0;rain_draw[24][50] = 0;rain_draw[25][50] = 0;rain_draw[26][50] = 0;rain_draw[27][50] = 0;rain_draw[28][50] = 0;rain_draw[29][50] = 0;rain_draw[30][50] = 0;rain_draw[31][50] = 0;rain_draw[32][50] = 0;rain_draw[33][50] = 0;rain_draw[34][50] = 0;rain_draw[35][50] = 0;rain_draw[36][50] = 0;rain_draw[37][50] = 1;rain_draw[38][50] = 1;rain_draw[39][50] = 1;rain_draw[40][50] = 0;rain_draw[41][50] = 0;rain_draw[42][50] = 0;rain_draw[43][50] = 0;rain_draw[44][50] = 0;rain_draw[45][50] = 0;rain_draw[46][50] = 0;rain_draw[47][50] = 0;rain_draw[48][50] = 0;rain_draw[49][50] = 0;rain_draw[50][50] = 0;rain_draw[51][50] = 0;rain_draw[52][50] = 0;rain_draw[53][50] = 0;rain_draw[54][50] = 0;rain_draw[55][50] = 0;rain_draw[56][50] = 0;rain_draw[57][50] = 0;rain_draw[58][50] = 0;rain_draw[59][50] = 0;rain_draw[60][50] = 0;rain_draw[61][50] = 0;rain_draw[62][50] = 0;rain_draw[63][50] = 1;rain_draw[64][50] = 1;rain_draw[65][50] = 1;rain_draw[66][50] = 0;rain_draw[67][50] = 0;rain_draw[68][50] = 0;rain_draw[69][50] = 0;rain_draw[70][50] = 0;rain_draw[71][50] = 0;rain_draw[72][50] = 0;rain_draw[73][50] = 0;rain_draw[74][50] = 0;rain_draw[75][50] = 0;rain_draw[76][50] = 0;rain_draw[77][50] = 0;rain_draw[78][50] = 0;rain_draw[79][50] = 0;rain_draw[80][50] = 0;rain_draw[81][50] = 0;rain_draw[82][50] = 0;rain_draw[83][50] = 0;rain_draw[84][50] = 0;rain_draw[85][50] = 0;rain_draw[86][50] = 0;rain_draw[87][50] = 0;rain_draw[88][50] = 0;rain_draw[89][50] = 0;rain_draw[90][50] = 0;rain_draw[91][50] = 0;rain_draw[92][50] = 0;rain_draw[93][50] = 0;rain_draw[94][50] = 0;rain_draw[95][50] = 0;
        rain_draw[0][51] = 0;rain_draw[1][51] = 0;rain_draw[2][51] = 0;rain_draw[3][51] = 0;rain_draw[4][51] = 0;rain_draw[5][51] = 0;rain_draw[6][51] = 0;rain_draw[7][51] = 0;rain_draw[8][51] = 0;rain_draw[9][51] = 0;rain_draw[10][51] = 0;rain_draw[11][51] = 0;rain_draw[12][51] = 0;rain_draw[13][51] = 0;rain_draw[14][51] = 0;rain_draw[15][51] = 0;rain_draw[16][51] = 0;rain_draw[17][51] = 0;rain_draw[18][51] = 0;rain_draw[19][51] = 0;rain_draw[20][51] = 0;rain_draw[21][51] = 0;rain_draw[22][51] = 0;rain_draw[23][51] = 0;rain_draw[24][51] = 0;rain_draw[25][51] = 0;rain_draw[26][51] = 0;rain_draw[27][51] = 0;rain_draw[28][51] = 0;rain_draw[29][51] = 0;rain_draw[30][51] = 0;rain_draw[31][51] = 0;rain_draw[32][51] = 0;rain_draw[33][51] = 0;rain_draw[34][51] = 0;rain_draw[35][51] = 0;rain_draw[36][51] = 1;rain_draw[37][51] = 1;rain_draw[38][51] = 1;rain_draw[39][51] = 0;rain_draw[40][51] = 0;rain_draw[41][51] = 0;rain_draw[42][51] = 0;rain_draw[43][51] = 0;rain_draw[44][51] = 0;rain_draw[45][51] = 0;rain_draw[46][51] = 0;rain_draw[47][51] = 0;rain_draw[48][51] = 0;rain_draw[49][51] = 0;rain_draw[50][51] = 0;rain_draw[51][51] = 0;rain_draw[52][51] = 0;rain_draw[53][51] = 0;rain_draw[54][51] = 0;rain_draw[55][51] = 0;rain_draw[56][51] = 0;rain_draw[57][51] = 0;rain_draw[58][51] = 0;rain_draw[59][51] = 0;rain_draw[60][51] = 0;rain_draw[61][51] = 0;rain_draw[62][51] = 1;rain_draw[63][51] = 1;rain_draw[64][51] = 1;rain_draw[65][51] = 0;rain_draw[66][51] = 0;rain_draw[67][51] = 0;rain_draw[68][51] = 0;rain_draw[69][51] = 0;rain_draw[70][51] = 0;rain_draw[71][51] = 0;rain_draw[72][51] = 0;rain_draw[73][51] = 0;rain_draw[74][51] = 0;rain_draw[75][51] = 0;rain_draw[76][51] = 0;rain_draw[77][51] = 0;rain_draw[78][51] = 0;rain_draw[79][51] = 0;rain_draw[80][51] = 0;rain_draw[81][51] = 0;rain_draw[82][51] = 0;rain_draw[83][51] = 0;rain_draw[84][51] = 0;rain_draw[85][51] = 0;rain_draw[86][51] = 0;rain_draw[87][51] = 0;rain_draw[88][51] = 0;rain_draw[89][51] = 0;rain_draw[90][51] = 0;rain_draw[91][51] = 0;rain_draw[92][51] = 0;rain_draw[93][51] = 0;rain_draw[94][51] = 0;rain_draw[95][51] = 0;
        rain_draw[0][52] = 0;rain_draw[1][52] = 0;rain_draw[2][52] = 0;rain_draw[3][52] = 0;rain_draw[4][52] = 0;rain_draw[5][52] = 0;rain_draw[6][52] = 0;rain_draw[7][52] = 0;rain_draw[8][52] = 0;rain_draw[9][52] = 0;rain_draw[10][52] = 0;rain_draw[11][52] = 0;rain_draw[12][52] = 0;rain_draw[13][52] = 0;rain_draw[14][52] = 0;rain_draw[15][52] = 0;rain_draw[16][52] = 0;rain_draw[17][52] = 0;rain_draw[18][52] = 0;rain_draw[19][52] = 0;rain_draw[20][52] = 0;rain_draw[21][52] = 0;rain_draw[22][52] = 0;rain_draw[23][52] = 0;rain_draw[24][52] = 0;rain_draw[25][52] = 0;rain_draw[26][52] = 0;rain_draw[27][52] = 0;rain_draw[28][52] = 0;rain_draw[29][52] = 0;rain_draw[30][52] = 0;rain_draw[31][52] = 0;rain_draw[32][52] = 0;rain_draw[33][52] = 0;rain_draw[34][52] = 0;rain_draw[35][52] = 1;rain_draw[36][52] = 1;rain_draw[37][52] = 1;rain_draw[38][52] = 0;rain_draw[39][52] = 0;rain_draw[40][52] = 0;rain_draw[41][52] = 0;rain_draw[42][52] = 0;rain_draw[43][52] = 0;rain_draw[44][52] = 0;rain_draw[45][52] = 0;rain_draw[46][52] = 0;rain_draw[47][52] = 0;rain_draw[48][52] = 0;rain_draw[49][52] = 0;rain_draw[50][52] = 0;rain_draw[51][52] = 0;rain_draw[52][52] = 0;rain_draw[53][52] = 0;rain_draw[54][52] = 0;rain_draw[55][52] = 0;rain_draw[56][52] = 0;rain_draw[57][52] = 0;rain_draw[58][52] = 0;rain_draw[59][52] = 0;rain_draw[60][52] = 0;rain_draw[61][52] = 1;rain_draw[62][52] = 1;rain_draw[63][52] = 1;rain_draw[64][52] = 0;rain_draw[65][52] = 0;rain_draw[66][52] = 0;rain_draw[67][52] = 0;rain_draw[68][52] = 0;rain_draw[69][52] = 0;rain_draw[70][52] = 0;rain_draw[71][52] = 0;rain_draw[72][52] = 0;rain_draw[73][52] = 0;rain_draw[74][52] = 0;rain_draw[75][52] = 0;rain_draw[76][52] = 0;rain_draw[77][52] = 0;rain_draw[78][52] = 0;rain_draw[79][52] = 0;rain_draw[80][52] = 0;rain_draw[81][52] = 0;rain_draw[82][52] = 0;rain_draw[83][52] = 0;rain_draw[84][52] = 0;rain_draw[85][52] = 0;rain_draw[86][52] = 0;rain_draw[87][52] = 0;rain_draw[88][52] = 0;rain_draw[89][52] = 0;rain_draw[90][52] = 0;rain_draw[91][52] = 0;rain_draw[92][52] = 0;rain_draw[93][52] = 0;rain_draw[94][52] = 0;rain_draw[95][52] = 0;
        rain_draw[0][53] = 0;rain_draw[1][53] = 0;rain_draw[2][53] = 0;rain_draw[3][53] = 0;rain_draw[4][53] = 0;rain_draw[5][53] = 0;rain_draw[6][53] = 0;rain_draw[7][53] = 0;rain_draw[8][53] = 0;rain_draw[9][53] = 0;rain_draw[10][53] = 0;rain_draw[11][53] = 0;rain_draw[12][53] = 0;rain_draw[13][53] = 0;rain_draw[14][53] = 0;rain_draw[15][53] = 0;rain_draw[16][53] = 0;rain_draw[17][53] = 0;rain_draw[18][53] = 0;rain_draw[19][53] = 0;rain_draw[20][53] = 0;rain_draw[21][53] = 0;rain_draw[22][53] = 0;rain_draw[23][53] = 0;rain_draw[24][53] = 0;rain_draw[25][53] = 0;rain_draw[26][53] = 0;rain_draw[27][53] = 0;rain_draw[28][53] = 0;rain_draw[29][53] = 0;rain_draw[30][53] = 0;rain_draw[31][53] = 0;rain_draw[32][53] = 0;rain_draw[33][53] = 0;rain_draw[34][53] = 0;rain_draw[35][53] = 0;rain_draw[36][53] = 0;rain_draw[37][53] = 0;rain_draw[38][53] = 0;rain_draw[39][53] = 0;rain_draw[40][53] = 0;rain_draw[41][53] = 0;rain_draw[42][53] = 0;rain_draw[43][53] = 0;rain_draw[44][53] = 0;rain_draw[45][53] = 0;rain_draw[46][53] = 0;rain_draw[47][53] = 0;rain_draw[48][53] = 0;rain_draw[49][53] = 0;rain_draw[50][53] = 0;rain_draw[51][53] = 0;rain_draw[52][53] = 0;rain_draw[53][53] = 0;rain_draw[54][53] = 0;rain_draw[55][53] = 0;rain_draw[56][53] = 0;rain_draw[57][53] = 0;rain_draw[58][53] = 0;rain_draw[59][53] = 0;rain_draw[60][53] = 1;rain_draw[61][53] = 1;rain_draw[62][53] = 1;rain_draw[63][53] = 0;rain_draw[64][53] = 0;rain_draw[65][53] = 0;rain_draw[66][53] = 0;rain_draw[67][53] = 0;rain_draw[68][53] = 0;rain_draw[69][53] = 0;rain_draw[70][53] = 0;rain_draw[71][53] = 0;rain_draw[72][53] = 0;rain_draw[73][53] = 0;rain_draw[74][53] = 0;rain_draw[75][53] = 0;rain_draw[76][53] = 0;rain_draw[77][53] = 0;rain_draw[78][53] = 0;rain_draw[79][53] = 0;rain_draw[80][53] = 0;rain_draw[81][53] = 0;rain_draw[82][53] = 0;rain_draw[83][53] = 0;rain_draw[84][53] = 0;rain_draw[85][53] = 0;rain_draw[86][53] = 0;rain_draw[87][53] = 0;rain_draw[88][53] = 0;rain_draw[89][53] = 0;rain_draw[90][53] = 0;rain_draw[91][53] = 0;rain_draw[92][53] = 0;rain_draw[93][53] = 0;rain_draw[94][53] = 0;rain_draw[95][53] = 0;
        rain_draw[0][54] = 0;rain_draw[1][54] = 0;rain_draw[2][54] = 0;rain_draw[3][54] = 0;rain_draw[4][54] = 0;rain_draw[5][54] = 0;rain_draw[6][54] = 0;rain_draw[7][54] = 0;rain_draw[8][54] = 0;rain_draw[9][54] = 0;rain_draw[10][54] = 0;rain_draw[11][54] = 0;rain_draw[12][54] = 0;rain_draw[13][54] = 0;rain_draw[14][54] = 0;rain_draw[15][54] = 0;rain_draw[16][54] = 0;rain_draw[17][54] = 0;rain_draw[18][54] = 0;rain_draw[19][54] = 0;rain_draw[20][54] = 0;rain_draw[21][54] = 0;rain_draw[22][54] = 0;rain_draw[23][54] = 0;rain_draw[24][54] = 0;rain_draw[25][54] = 0;rain_draw[26][54] = 0;rain_draw[27][54] = 0;rain_draw[28][54] = 0;rain_draw[29][54] = 0;rain_draw[30][54] = 0;rain_draw[31][54] = 0;rain_draw[32][54] = 0;rain_draw[33][54] = 0;rain_draw[34][54] = 0;rain_draw[35][54] = 0;rain_draw[36][54] = 0;rain_draw[37][54] = 0;rain_draw[38][54] = 0;rain_draw[39][54] = 0;rain_draw[40][54] = 0;rain_draw[41][54] = 0;rain_draw[42][54] = 0;rain_draw[43][54] = 0;rain_draw[44][54] = 0;rain_draw[45][54] = 0;rain_draw[46][54] = 0;rain_draw[47][54] = 0;rain_draw[48][54] = 0;rain_draw[49][54] = 0;rain_draw[50][54] = 0;rain_draw[51][54] = 0;rain_draw[52][54] = 0;rain_draw[53][54] = 0;rain_draw[54][54] = 0;rain_draw[55][54] = 0;rain_draw[56][54] = 0;rain_draw[57][54] = 0;rain_draw[58][54] = 0;rain_draw[59][54] = 1;rain_draw[60][54] = 1;rain_draw[61][54] = 1;rain_draw[62][54] = 0;rain_draw[63][54] = 0;rain_draw[64][54] = 0;rain_draw[65][54] = 0;rain_draw[66][54] = 0;rain_draw[67][54] = 0;rain_draw[68][54] = 0;rain_draw[69][54] = 0;rain_draw[70][54] = 0;rain_draw[71][54] = 0;rain_draw[72][54] = 0;rain_draw[73][54] = 0;rain_draw[74][54] = 0;rain_draw[75][54] = 0;rain_draw[76][54] = 0;rain_draw[77][54] = 0;rain_draw[78][54] = 0;rain_draw[79][54] = 0;rain_draw[80][54] = 0;rain_draw[81][54] = 0;rain_draw[82][54] = 0;rain_draw[83][54] = 0;rain_draw[84][54] = 0;rain_draw[85][54] = 0;rain_draw[86][54] = 0;rain_draw[87][54] = 0;rain_draw[88][54] = 0;rain_draw[89][54] = 0;rain_draw[90][54] = 0;rain_draw[91][54] = 0;rain_draw[92][54] = 0;rain_draw[93][54] = 0;rain_draw[94][54] = 0;rain_draw[95][54] = 0;
        rain_draw[0][55] = 0;rain_draw[1][55] = 0;rain_draw[2][55] = 0;rain_draw[3][55] = 0;rain_draw[4][55] = 0;rain_draw[5][55] = 0;rain_draw[6][55] = 0;rain_draw[7][55] = 0;rain_draw[8][55] = 0;rain_draw[9][55] = 0;rain_draw[10][55] = 0;rain_draw[11][55] = 0;rain_draw[12][55] = 0;rain_draw[13][55] = 0;rain_draw[14][55] = 0;rain_draw[15][55] = 0;rain_draw[16][55] = 0;rain_draw[17][55] = 0;rain_draw[18][55] = 0;rain_draw[19][55] = 0;rain_draw[20][55] = 0;rain_draw[21][55] = 0;rain_draw[22][55] = 0;rain_draw[23][55] = 0;rain_draw[24][55] = 0;rain_draw[25][55] = 0;rain_draw[26][55] = 0;rain_draw[27][55] = 0;rain_draw[28][55] = 0;rain_draw[29][55] = 0;rain_draw[30][55] = 0;rain_draw[31][55] = 0;rain_draw[32][55] = 0;rain_draw[33][55] = 0;rain_draw[34][55] = 0;rain_draw[35][55] = 0;rain_draw[36][55] = 0;rain_draw[37][55] = 0;rain_draw[38][55] = 0;rain_draw[39][55] = 0;rain_draw[40][55] = 0;rain_draw[41][55] = 0;rain_draw[42][55] = 0;rain_draw[43][55] = 0;rain_draw[44][55] = 0;rain_draw[45][55] = 0;rain_draw[46][55] = 0;rain_draw[47][55] = 0;rain_draw[48][55] = 0;rain_draw[49][55] = 0;rain_draw[50][55] = 0;rain_draw[51][55] = 0;rain_draw[52][55] = 0;rain_draw[53][55] = 0;rain_draw[54][55] = 0;rain_draw[55][55] = 0;rain_draw[56][55] = 0;rain_draw[57][55] = 0;rain_draw[58][55] = 1;rain_draw[59][55] = 1;rain_draw[60][55] = 1;rain_draw[61][55] = 0;rain_draw[62][55] = 0;rain_draw[63][55] = 0;rain_draw[64][55] = 0;rain_draw[65][55] = 0;rain_draw[66][55] = 0;rain_draw[67][55] = 0;rain_draw[68][55] = 0;rain_draw[69][55] = 0;rain_draw[70][55] = 0;rain_draw[71][55] = 0;rain_draw[72][55] = 0;rain_draw[73][55] = 0;rain_draw[74][55] = 0;rain_draw[75][55] = 0;rain_draw[76][55] = 0;rain_draw[77][55] = 0;rain_draw[78][55] = 0;rain_draw[79][55] = 0;rain_draw[80][55] = 0;rain_draw[81][55] = 1;rain_draw[82][55] = 1;rain_draw[83][55] = 1;rain_draw[84][55] = 0;rain_draw[85][55] = 0;rain_draw[86][55] = 0;rain_draw[87][55] = 0;rain_draw[88][55] = 0;rain_draw[89][55] = 0;rain_draw[90][55] = 0;rain_draw[91][55] = 0;rain_draw[92][55] = 0;rain_draw[93][55] = 0;rain_draw[94][55] = 0;rain_draw[95][55] = 0;
        rain_draw[0][56] = 0;rain_draw[1][56] = 0;rain_draw[2][56] = 0;rain_draw[3][56] = 0;rain_draw[4][56] = 0;rain_draw[5][56] = 0;rain_draw[6][56] = 0;rain_draw[7][56] = 0;rain_draw[8][56] = 0;rain_draw[9][56] = 0;rain_draw[10][56] = 0;rain_draw[11][56] = 0;rain_draw[12][56] = 0;rain_draw[13][56] = 0;rain_draw[14][56] = 0;rain_draw[15][56] = 0;rain_draw[16][56] = 0;rain_draw[17][56] = 0;rain_draw[18][56] = 0;rain_draw[19][56] = 0;rain_draw[20][56] = 0;rain_draw[21][56] = 0;rain_draw[22][56] = 0;rain_draw[23][56] = 0;rain_draw[24][56] = 0;rain_draw[25][56] = 0;rain_draw[26][56] = 0;rain_draw[27][56] = 0;rain_draw[28][56] = 0;rain_draw[29][56] = 0;rain_draw[30][56] = 0;rain_draw[31][56] = 0;rain_draw[32][56] = 0;rain_draw[33][56] = 0;rain_draw[34][56] = 0;rain_draw[35][56] = 0;rain_draw[36][56] = 0;rain_draw[37][56] = 0;rain_draw[38][56] = 0;rain_draw[39][56] = 0;rain_draw[40][56] = 0;rain_draw[41][56] = 0;rain_draw[42][56] = 0;rain_draw[43][56] = 0;rain_draw[44][56] = 0;rain_draw[45][56] = 0;rain_draw[46][56] = 0;rain_draw[47][56] = 0;rain_draw[48][56] = 0;rain_draw[49][56] = 0;rain_draw[50][56] = 0;rain_draw[51][56] = 0;rain_draw[52][56] = 0;rain_draw[53][56] = 0;rain_draw[54][56] = 0;rain_draw[55][56] = 0;rain_draw[56][56] = 0;rain_draw[57][56] = 1;rain_draw[58][56] = 1;rain_draw[59][56] = 1;rain_draw[60][56] = 0;rain_draw[61][56] = 0;rain_draw[62][56] = 0;rain_draw[63][56] = 0;rain_draw[64][56] = 0;rain_draw[65][56] = 0;rain_draw[66][56] = 0;rain_draw[67][56] = 0;rain_draw[68][56] = 0;rain_draw[69][56] = 0;rain_draw[70][56] = 0;rain_draw[71][56] = 0;rain_draw[72][56] = 0;rain_draw[73][56] = 0;rain_draw[74][56] = 0;rain_draw[75][56] = 0;rain_draw[76][56] = 0;rain_draw[77][56] = 0;rain_draw[78][56] = 0;rain_draw[79][56] = 0;rain_draw[80][56] = 1;rain_draw[81][56] = 1;rain_draw[82][56] = 1;rain_draw[83][56] = 0;rain_draw[84][56] = 0;rain_draw[85][56] = 0;rain_draw[86][56] = 0;rain_draw[87][56] = 0;rain_draw[88][56] = 0;rain_draw[89][56] = 0;rain_draw[90][56] = 0;rain_draw[91][56] = 0;rain_draw[92][56] = 0;rain_draw[93][56] = 0;rain_draw[94][56] = 0;rain_draw[95][56] = 0;
        rain_draw[0][57] = 0;rain_draw[1][57] = 0;rain_draw[2][57] = 0;rain_draw[3][57] = 0;rain_draw[4][57] = 0;rain_draw[5][57] = 0;rain_draw[6][57] = 0;rain_draw[7][57] = 0;rain_draw[8][57] = 0;rain_draw[9][57] = 0;rain_draw[10][57] = 0;rain_draw[11][57] = 0;rain_draw[12][57] = 0;rain_draw[13][57] = 0;rain_draw[14][57] = 0;rain_draw[15][57] = 0;rain_draw[16][57] = 0;rain_draw[17][57] = 0;rain_draw[18][57] = 0;rain_draw[19][57] = 0;rain_draw[20][57] = 0;rain_draw[21][57] = 0;rain_draw[22][57] = 0;rain_draw[23][57] = 0;rain_draw[24][57] = 0;rain_draw[25][57] = 0;rain_draw[26][57] = 0;rain_draw[27][57] = 0;rain_draw[28][57] = 0;rain_draw[29][57] = 0;rain_draw[30][57] = 0;rain_draw[31][57] = 0;rain_draw[32][57] = 0;rain_draw[33][57] = 0;rain_draw[34][57] = 0;rain_draw[35][57] = 0;rain_draw[36][57] = 0;rain_draw[37][57] = 0;rain_draw[38][57] = 0;rain_draw[39][57] = 0;rain_draw[40][57] = 0;rain_draw[41][57] = 0;rain_draw[42][57] = 0;rain_draw[43][57] = 0;rain_draw[44][57] = 0;rain_draw[45][57] = 0;rain_draw[46][57] = 0;rain_draw[47][57] = 0;rain_draw[48][57] = 0;rain_draw[49][57] = 0;rain_draw[50][57] = 0;rain_draw[51][57] = 0;rain_draw[52][57] = 0;rain_draw[53][57] = 0;rain_draw[54][57] = 0;rain_draw[55][57] = 0;rain_draw[56][57] = 0;rain_draw[57][57] = 0;rain_draw[58][57] = 0;rain_draw[59][57] = 0;rain_draw[60][57] = 0;rain_draw[61][57] = 0;rain_draw[62][57] = 0;rain_draw[63][57] = 0;rain_draw[64][57] = 0;rain_draw[65][57] = 0;rain_draw[66][57] = 0;rain_draw[67][57] = 0;rain_draw[68][57] = 0;rain_draw[69][57] = 0;rain_draw[70][57] = 0;rain_draw[71][57] = 0;rain_draw[72][57] = 0;rain_draw[73][57] = 0;rain_draw[74][57] = 0;rain_draw[75][57] = 0;rain_draw[76][57] = 0;rain_draw[77][57] = 0;rain_draw[78][57] = 0;rain_draw[79][57] = 1;rain_draw[80][57] = 1;rain_draw[81][57] = 1;rain_draw[82][57] = 0;rain_draw[83][57] = 0;rain_draw[84][57] = 0;rain_draw[85][57] = 0;rain_draw[86][57] = 0;rain_draw[87][57] = 0;rain_draw[88][57] = 0;rain_draw[89][57] = 0;rain_draw[90][57] = 0;rain_draw[91][57] = 0;rain_draw[92][57] = 0;rain_draw[93][57] = 0;rain_draw[94][57] = 0;rain_draw[95][57] = 0;
        rain_draw[0][58] = 0;rain_draw[1][58] = 0;rain_draw[2][58] = 0;rain_draw[3][58] = 0;rain_draw[4][58] = 0;rain_draw[5][58] = 0;rain_draw[6][58] = 0;rain_draw[7][58] = 0;rain_draw[8][58] = 0;rain_draw[9][58] = 0;rain_draw[10][58] = 0;rain_draw[11][58] = 0;rain_draw[12][58] = 0;rain_draw[13][58] = 0;rain_draw[14][58] = 0;rain_draw[15][58] = 0;rain_draw[16][58] = 0;rain_draw[17][58] = 0;rain_draw[18][58] = 0;rain_draw[19][58] = 0;rain_draw[20][58] = 0;rain_draw[21][58] = 0;rain_draw[22][58] = 0;rain_draw[23][58] = 0;rain_draw[24][58] = 0;rain_draw[25][58] = 0;rain_draw[26][58] = 0;rain_draw[27][58] = 0;rain_draw[28][58] = 0;rain_draw[29][58] = 0;rain_draw[30][58] = 0;rain_draw[31][58] = 0;rain_draw[32][58] = 0;rain_draw[33][58] = 0;rain_draw[34][58] = 0;rain_draw[35][58] = 0;rain_draw[36][58] = 0;rain_draw[37][58] = 0;rain_draw[38][58] = 0;rain_draw[39][58] = 0;rain_draw[40][58] = 0;rain_draw[41][58] = 0;rain_draw[42][58] = 0;rain_draw[43][58] = 0;rain_draw[44][58] = 0;rain_draw[45][58] = 0;rain_draw[46][58] = 0;rain_draw[47][58] = 0;rain_draw[48][58] = 0;rain_draw[49][58] = 0;rain_draw[50][58] = 0;rain_draw[51][58] = 0;rain_draw[52][58] = 0;rain_draw[53][58] = 0;rain_draw[54][58] = 0;rain_draw[55][58] = 0;rain_draw[56][58] = 0;rain_draw[57][58] = 0;rain_draw[58][58] = 0;rain_draw[59][58] = 0;rain_draw[60][58] = 0;rain_draw[61][58] = 0;rain_draw[62][58] = 0;rain_draw[63][58] = 0;rain_draw[64][58] = 0;rain_draw[65][58] = 0;rain_draw[66][58] = 0;rain_draw[67][58] = 0;rain_draw[68][58] = 0;rain_draw[69][58] = 0;rain_draw[70][58] = 0;rain_draw[71][58] = 0;rain_draw[72][58] = 0;rain_draw[73][58] = 0;rain_draw[74][58] = 0;rain_draw[75][58] = 0;rain_draw[76][58] = 0;rain_draw[77][58] = 0;rain_draw[78][58] = 1;rain_draw[79][58] = 1;rain_draw[80][58] = 1;rain_draw[81][58] = 0;rain_draw[82][58] = 0;rain_draw[83][58] = 0;rain_draw[84][58] = 0;rain_draw[85][58] = 0;rain_draw[86][58] = 0;rain_draw[87][58] = 0;rain_draw[88][58] = 0;rain_draw[89][58] = 0;rain_draw[90][58] = 0;rain_draw[91][58] = 0;rain_draw[92][58] = 0;rain_draw[93][58] = 0;rain_draw[94][58] = 0;rain_draw[95][58] = 0;
        rain_draw[0][59] = 0;rain_draw[1][59] = 0;rain_draw[2][59] = 0;rain_draw[3][59] = 0;rain_draw[4][59] = 0;rain_draw[5][59] = 0;rain_draw[6][59] = 0;rain_draw[7][59] = 0;rain_draw[8][59] = 0;rain_draw[9][59] = 0;rain_draw[10][59] = 0;rain_draw[11][59] = 0;rain_draw[12][59] = 0;rain_draw[13][59] = 0;rain_draw[14][59] = 0;rain_draw[15][59] = 0;rain_draw[16][59] = 0;rain_draw[17][59] = 0;rain_draw[18][59] = 0;rain_draw[19][59] = 0;rain_draw[20][59] = 0;rain_draw[21][59] = 0;rain_draw[22][59] = 0;rain_draw[23][59] = 0;rain_draw[24][59] = 0;rain_draw[25][59] = 0;rain_draw[26][59] = 0;rain_draw[27][59] = 0;rain_draw[28][59] = 0;rain_draw[29][59] = 0;rain_draw[30][59] = 0;rain_draw[31][59] = 0;rain_draw[32][59] = 0;rain_draw[33][59] = 0;rain_draw[34][59] = 0;rain_draw[35][59] = 0;rain_draw[36][59] = 0;rain_draw[37][59] = 0;rain_draw[38][59] = 0;rain_draw[39][59] = 0;rain_draw[40][59] = 0;rain_draw[41][59] = 0;rain_draw[42][59] = 0;rain_draw[43][59] = 0;rain_draw[44][59] = 0;rain_draw[45][59] = 0;rain_draw[46][59] = 0;rain_draw[47][59] = 0;rain_draw[48][59] = 0;rain_draw[49][59] = 0;rain_draw[50][59] = 0;rain_draw[51][59] = 0;rain_draw[52][59] = 0;rain_draw[53][59] = 0;rain_draw[54][59] = 0;rain_draw[55][59] = 0;rain_draw[56][59] = 0;rain_draw[57][59] = 0;rain_draw[58][59] = 0;rain_draw[59][59] = 0;rain_draw[60][59] = 0;rain_draw[61][59] = 0;rain_draw[62][59] = 0;rain_draw[63][59] = 0;rain_draw[64][59] = 0;rain_draw[65][59] = 0;rain_draw[66][59] = 0;rain_draw[67][59] = 0;rain_draw[68][59] = 0;rain_draw[69][59] = 0;rain_draw[70][59] = 0;rain_draw[71][59] = 0;rain_draw[72][59] = 0;rain_draw[73][59] = 0;rain_draw[74][59] = 0;rain_draw[75][59] = 0;rain_draw[76][59] = 0;rain_draw[77][59] = 1;rain_draw[78][59] = 1;rain_draw[79][59] = 1;rain_draw[80][59] = 0;rain_draw[81][59] = 0;rain_draw[82][59] = 0;rain_draw[83][59] = 0;rain_draw[84][59] = 0;rain_draw[85][59] = 0;rain_draw[86][59] = 0;rain_draw[87][59] = 0;rain_draw[88][59] = 0;rain_draw[89][59] = 0;rain_draw[90][59] = 0;rain_draw[91][59] = 0;rain_draw[92][59] = 0;rain_draw[93][59] = 0;rain_draw[94][59] = 0;rain_draw[95][59] = 0;
        rain_draw[0][60] = 0;rain_draw[1][60] = 0;rain_draw[2][60] = 0;rain_draw[3][60] = 0;rain_draw[4][60] = 0;rain_draw[5][60] = 0;rain_draw[6][60] = 0;rain_draw[7][60] = 0;rain_draw[8][60] = 0;rain_draw[9][60] = 0;rain_draw[10][60] = 0;rain_draw[11][60] = 0;rain_draw[12][60] = 0;rain_draw[13][60] = 0;rain_draw[14][60] = 0;rain_draw[15][60] = 0;rain_draw[16][60] = 0;rain_draw[17][60] = 0;rain_draw[18][60] = 0;rain_draw[19][60] = 0;rain_draw[20][60] = 0;rain_draw[21][60] = 0;rain_draw[22][60] = 0;rain_draw[23][60] = 0;rain_draw[24][60] = 0;rain_draw[25][60] = 0;rain_draw[26][60] = 0;rain_draw[27][60] = 0;rain_draw[28][60] = 0;rain_draw[29][60] = 0;rain_draw[30][60] = 0;rain_draw[31][60] = 0;rain_draw[32][60] = 0;rain_draw[33][60] = 0;rain_draw[34][60] = 0;rain_draw[35][60] = 0;rain_draw[36][60] = 0;rain_draw[37][60] = 0;rain_draw[38][60] = 0;rain_draw[39][60] = 0;rain_draw[40][60] = 0;rain_draw[41][60] = 0;rain_draw[42][60] = 0;rain_draw[43][60] = 0;rain_draw[44][60] = 0;rain_draw[45][60] = 0;rain_draw[46][60] = 0;rain_draw[47][60] = 0;rain_draw[48][60] = 0;rain_draw[49][60] = 0;rain_draw[50][60] = 0;rain_draw[51][60] = 0;rain_draw[52][60] = 0;rain_draw[53][60] = 0;rain_draw[54][60] = 0;rain_draw[55][60] = 0;rain_draw[56][60] = 0;rain_draw[57][60] = 0;rain_draw[58][60] = 0;rain_draw[59][60] = 0;rain_draw[60][60] = 0;rain_draw[61][60] = 0;rain_draw[62][60] = 0;rain_draw[63][60] = 0;rain_draw[64][60] = 0;rain_draw[65][60] = 0;rain_draw[66][60] = 0;rain_draw[67][60] = 0;rain_draw[68][60] = 0;rain_draw[69][60] = 0;rain_draw[70][60] = 0;rain_draw[71][60] = 0;rain_draw[72][60] = 0;rain_draw[73][60] = 0;rain_draw[74][60] = 0;rain_draw[75][60] = 0;rain_draw[76][60] = 1;rain_draw[77][60] = 1;rain_draw[78][60] = 1;rain_draw[79][60] = 0;rain_draw[80][60] = 0;rain_draw[81][60] = 0;rain_draw[82][60] = 0;rain_draw[83][60] = 0;rain_draw[84][60] = 0;rain_draw[85][60] = 0;rain_draw[86][60] = 0;rain_draw[87][60] = 0;rain_draw[88][60] = 0;rain_draw[89][60] = 0;rain_draw[90][60] = 0;rain_draw[91][60] = 0;rain_draw[92][60] = 0;rain_draw[93][60] = 0;rain_draw[94][60] = 0;rain_draw[95][60] = 0;
        rain_draw[0][61] = 0;rain_draw[1][61] = 0;rain_draw[2][61] = 0;rain_draw[3][61] = 0;rain_draw[4][61] = 0;rain_draw[5][61] = 0;rain_draw[6][61] = 0;rain_draw[7][61] = 0;rain_draw[8][61] = 0;rain_draw[9][61] = 0;rain_draw[10][61] = 0;rain_draw[11][61] = 0;rain_draw[12][61] = 0;rain_draw[13][61] = 0;rain_draw[14][61] = 0;rain_draw[15][61] = 0;rain_draw[16][61] = 0;rain_draw[17][61] = 0;rain_draw[18][61] = 0;rain_draw[19][61] = 0;rain_draw[20][61] = 0;rain_draw[21][61] = 0;rain_draw[22][61] = 0;rain_draw[23][61] = 0;rain_draw[24][61] = 0;rain_draw[25][61] = 0;rain_draw[26][61] = 0;rain_draw[27][61] = 0;rain_draw[28][61] = 0;rain_draw[29][61] = 0;rain_draw[30][61] = 0;rain_draw[31][61] = 0;rain_draw[32][61] = 0;rain_draw[33][61] = 0;rain_draw[34][61] = 0;rain_draw[35][61] = 0;rain_draw[36][61] = 0;rain_draw[37][61] = 0;rain_draw[38][61] = 0;rain_draw[39][61] = 0;rain_draw[40][61] = 0;rain_draw[41][61] = 0;rain_draw[42][61] = 0;rain_draw[43][61] = 0;rain_draw[44][61] = 0;rain_draw[45][61] = 0;rain_draw[46][61] = 0;rain_draw[47][61] = 0;rain_draw[48][61] = 0;rain_draw[49][61] = 0;rain_draw[50][61] = 0;rain_draw[51][61] = 0;rain_draw[52][61] = 0;rain_draw[53][61] = 0;rain_draw[54][61] = 0;rain_draw[55][61] = 0;rain_draw[56][61] = 0;rain_draw[57][61] = 0;rain_draw[58][61] = 0;rain_draw[59][61] = 0;rain_draw[60][61] = 0;rain_draw[61][61] = 0;rain_draw[62][61] = 0;rain_draw[63][61] = 0;rain_draw[64][61] = 0;rain_draw[65][61] = 0;rain_draw[66][61] = 0;rain_draw[67][61] = 0;rain_draw[68][61] = 0;rain_draw[69][61] = 0;rain_draw[70][61] = 0;rain_draw[71][61] = 0;rain_draw[72][61] = 0;rain_draw[73][61] = 0;rain_draw[74][61] = 0;rain_draw[75][61] = 1;rain_draw[76][61] = 1;rain_draw[77][61] = 1;rain_draw[78][61] = 0;rain_draw[79][61] = 0;rain_draw[80][61] = 0;rain_draw[81][61] = 0;rain_draw[82][61] = 0;rain_draw[83][61] = 0;rain_draw[84][61] = 0;rain_draw[85][61] = 0;rain_draw[86][61] = 0;rain_draw[87][61] = 0;rain_draw[88][61] = 0;rain_draw[89][61] = 0;rain_draw[90][61] = 0;rain_draw[91][61] = 0;rain_draw[92][61] = 0;rain_draw[93][61] = 0;rain_draw[94][61] = 0;rain_draw[95][61] = 0;
        rain_draw[0][62] = 0;rain_draw[1][62] = 0;rain_draw[2][62] = 0;rain_draw[3][62] = 0;rain_draw[4][62] = 0;rain_draw[5][62] = 0;rain_draw[6][62] = 0;rain_draw[7][62] = 0;rain_draw[8][62] = 0;rain_draw[9][62] = 0;rain_draw[10][62] = 0;rain_draw[11][62] = 0;rain_draw[12][62] = 0;rain_draw[13][62] = 0;rain_draw[14][62] = 0;rain_draw[15][62] = 0;rain_draw[16][62] = 0;rain_draw[17][62] = 0;rain_draw[18][62] = 0;rain_draw[19][62] = 0;rain_draw[20][62] = 0;rain_draw[21][62] = 0;rain_draw[22][62] = 0;rain_draw[23][62] = 0;rain_draw[24][62] = 0;rain_draw[25][62] = 0;rain_draw[26][62] = 0;rain_draw[27][62] = 0;rain_draw[28][62] = 0;rain_draw[29][62] = 0;rain_draw[30][62] = 0;rain_draw[31][62] = 0;rain_draw[32][62] = 0;rain_draw[33][62] = 0;rain_draw[34][62] = 0;rain_draw[35][62] = 0;rain_draw[36][62] = 0;rain_draw[37][62] = 0;rain_draw[38][62] = 0;rain_draw[39][62] = 0;rain_draw[40][62] = 0;rain_draw[41][62] = 0;rain_draw[42][62] = 0;rain_draw[43][62] = 0;rain_draw[44][62] = 0;rain_draw[45][62] = 0;rain_draw[46][62] = 0;rain_draw[47][62] = 0;rain_draw[48][62] = 0;rain_draw[49][62] = 0;rain_draw[50][62] = 0;rain_draw[51][62] = 0;rain_draw[52][62] = 0;rain_draw[53][62] = 0;rain_draw[54][62] = 0;rain_draw[55][62] = 0;rain_draw[56][62] = 0;rain_draw[57][62] = 0;rain_draw[58][62] = 0;rain_draw[59][62] = 0;rain_draw[60][62] = 0;rain_draw[61][62] = 0;rain_draw[62][62] = 0;rain_draw[63][62] = 0;rain_draw[64][62] = 0;rain_draw[65][62] = 0;rain_draw[66][62] = 0;rain_draw[67][62] = 0;rain_draw[68][62] = 0;rain_draw[69][62] = 0;rain_draw[70][62] = 0;rain_draw[71][62] = 0;rain_draw[72][62] = 0;rain_draw[73][62] = 0;rain_draw[74][62] = 0;rain_draw[75][62] = 0;rain_draw[76][62] = 0;rain_draw[77][62] = 0;rain_draw[78][62] = 0;rain_draw[79][62] = 0;rain_draw[80][62] = 0;rain_draw[81][62] = 0;rain_draw[82][62] = 0;rain_draw[83][62] = 0;rain_draw[84][62] = 0;rain_draw[85][62] = 0;rain_draw[86][62] = 0;rain_draw[87][62] = 0;rain_draw[88][62] = 0;rain_draw[89][62] = 0;rain_draw[90][62] = 0;rain_draw[91][62] = 0;rain_draw[92][62] = 0;rain_draw[93][62] = 0;rain_draw[94][62] = 0;rain_draw[95][62] = 0;
        rain_draw[0][63] = 0;rain_draw[1][63] = 0;rain_draw[2][63] = 0;rain_draw[3][63] = 0;rain_draw[4][63] = 0;rain_draw[5][63] = 0;rain_draw[6][63] = 0;rain_draw[7][63] = 0;rain_draw[8][63] = 0;rain_draw[9][63] = 0;rain_draw[10][63] = 0;rain_draw[11][63] = 0;rain_draw[12][63] = 0;rain_draw[13][63] = 0;rain_draw[14][63] = 0;rain_draw[15][63] = 0;rain_draw[16][63] = 0;rain_draw[17][63] = 0;rain_draw[18][63] = 0;rain_draw[19][63] = 0;rain_draw[20][63] = 0;rain_draw[21][63] = 0;rain_draw[22][63] = 0;rain_draw[23][63] = 0;rain_draw[24][63] = 0;rain_draw[25][63] = 0;rain_draw[26][63] = 0;rain_draw[27][63] = 0;rain_draw[28][63] = 0;rain_draw[29][63] = 0;rain_draw[30][63] = 0;rain_draw[31][63] = 0;rain_draw[32][63] = 0;rain_draw[33][63] = 0;rain_draw[34][63] = 0;rain_draw[35][63] = 0;rain_draw[36][63] = 0;rain_draw[37][63] = 0;rain_draw[38][63] = 0;rain_draw[39][63] = 0;rain_draw[40][63] = 0;rain_draw[41][63] = 0;rain_draw[42][63] = 0;rain_draw[43][63] = 0;rain_draw[44][63] = 0;rain_draw[45][63] = 0;rain_draw[46][63] = 0;rain_draw[47][63] = 0;rain_draw[48][63] = 0;rain_draw[49][63] = 0;rain_draw[50][63] = 0;rain_draw[51][63] = 0;rain_draw[52][63] = 0;rain_draw[53][63] = 0;rain_draw[54][63] = 0;rain_draw[55][63] = 0;rain_draw[56][63] = 0;rain_draw[57][63] = 0;rain_draw[58][63] = 0;rain_draw[59][63] = 0;rain_draw[60][63] = 0;rain_draw[61][63] = 0;rain_draw[62][63] = 0;rain_draw[63][63] = 0;rain_draw[64][63] = 0;rain_draw[65][63] = 0;rain_draw[66][63] = 0;rain_draw[67][63] = 0;rain_draw[68][63] = 0;rain_draw[69][63] = 0;rain_draw[70][63] = 0;rain_draw[71][63] = 0;rain_draw[72][63] = 0;rain_draw[73][63] = 0;rain_draw[74][63] = 0;rain_draw[75][63] = 0;rain_draw[76][63] = 0;rain_draw[77][63] = 0;rain_draw[78][63] = 0;rain_draw[79][63] = 0;rain_draw[80][63] = 0;rain_draw[81][63] = 0;rain_draw[82][63] = 0;rain_draw[83][63] = 0;rain_draw[84][63] = 0;rain_draw[85][63] = 0;rain_draw[86][63] = 0;rain_draw[87][63] = 0;rain_draw[88][63] = 0;rain_draw[89][63] = 0;rain_draw[90][63] = 0;rain_draw[91][63] = 0;rain_draw[92][63] = 0;rain_draw[93][63] = 0;rain_draw[94][63] = 0;rain_draw[95][63] = 0;
        rain_draw[0][64] = 0;rain_draw[1][64] = 0;rain_draw[2][64] = 0;rain_draw[3][64] = 0;rain_draw[4][64] = 0;rain_draw[5][64] = 0;rain_draw[6][64] = 0;rain_draw[7][64] = 0;rain_draw[8][64] = 0;rain_draw[9][64] = 0;rain_draw[10][64] = 0;rain_draw[11][64] = 0;rain_draw[12][64] = 0;rain_draw[13][64] = 0;rain_draw[14][64] = 0;rain_draw[15][64] = 0;rain_draw[16][64] = 0;rain_draw[17][64] = 0;rain_draw[18][64] = 0;rain_draw[19][64] = 0;rain_draw[20][64] = 0;rain_draw[21][64] = 0;rain_draw[22][64] = 0;rain_draw[23][64] = 0;rain_draw[24][64] = 0;rain_draw[25][64] = 0;rain_draw[26][64] = 0;rain_draw[27][64] = 0;rain_draw[28][64] = 0;rain_draw[29][64] = 0;rain_draw[30][64] = 0;rain_draw[31][64] = 0;rain_draw[32][64] = 0;rain_draw[33][64] = 0;rain_draw[34][64] = 0;rain_draw[35][64] = 0;rain_draw[36][64] = 0;rain_draw[37][64] = 0;rain_draw[38][64] = 0;rain_draw[39][64] = 0;rain_draw[40][64] = 0;rain_draw[41][64] = 0;rain_draw[42][64] = 0;rain_draw[43][64] = 0;rain_draw[44][64] = 0;rain_draw[45][64] = 0;rain_draw[46][64] = 0;rain_draw[47][64] = 0;rain_draw[48][64] = 0;rain_draw[49][64] = 0;rain_draw[50][64] = 0;rain_draw[51][64] = 0;rain_draw[52][64] = 0;rain_draw[53][64] = 0;rain_draw[54][64] = 0;rain_draw[55][64] = 0;rain_draw[56][64] = 0;rain_draw[57][64] = 0;rain_draw[58][64] = 0;rain_draw[59][64] = 0;rain_draw[60][64] = 0;rain_draw[61][64] = 0;rain_draw[62][64] = 0;rain_draw[63][64] = 0;rain_draw[64][64] = 0;rain_draw[65][64] = 0;rain_draw[66][64] = 0;rain_draw[67][64] = 0;rain_draw[68][64] = 0;rain_draw[69][64] = 0;rain_draw[70][64] = 0;rain_draw[71][64] = 0;rain_draw[72][64] = 0;rain_draw[73][64] = 0;rain_draw[74][64] = 0;rain_draw[75][64] = 0;rain_draw[76][64] = 0;rain_draw[77][64] = 0;rain_draw[78][64] = 0;rain_draw[79][64] = 0;rain_draw[80][64] = 0;rain_draw[81][64] = 0;rain_draw[82][64] = 0;rain_draw[83][64] = 0;rain_draw[84][64] = 0;rain_draw[85][64] = 0;rain_draw[86][64] = 0;rain_draw[87][64] = 0;rain_draw[88][64] = 0;rain_draw[89][64] = 0;rain_draw[90][64] = 0;rain_draw[91][64] = 0;rain_draw[92][64] = 0;rain_draw[93][64] = 0;rain_draw[94][64] = 0;rain_draw[95][64] = 0;
        rain_draw[0][65] = 0;rain_draw[1][65] = 0;rain_draw[2][65] = 0;rain_draw[3][65] = 0;rain_draw[4][65] = 0;rain_draw[5][65] = 0;rain_draw[6][65] = 0;rain_draw[7][65] = 0;rain_draw[8][65] = 0;rain_draw[9][65] = 0;rain_draw[10][65] = 0;rain_draw[11][65] = 0;rain_draw[12][65] = 0;rain_draw[13][65] = 0;rain_draw[14][65] = 0;rain_draw[15][65] = 0;rain_draw[16][65] = 0;rain_draw[17][65] = 0;rain_draw[18][65] = 0;rain_draw[19][65] = 0;rain_draw[20][65] = 0;rain_draw[21][65] = 0;rain_draw[22][65] = 0;rain_draw[23][65] = 0;rain_draw[24][65] = 0;rain_draw[25][65] = 0;rain_draw[26][65] = 0;rain_draw[27][65] = 0;rain_draw[28][65] = 0;rain_draw[29][65] = 0;rain_draw[30][65] = 0;rain_draw[31][65] = 0;rain_draw[32][65] = 0;rain_draw[33][65] = 0;rain_draw[34][65] = 0;rain_draw[35][65] = 0;rain_draw[36][65] = 0;rain_draw[37][65] = 0;rain_draw[38][65] = 0;rain_draw[39][65] = 0;rain_draw[40][65] = 0;rain_draw[41][65] = 0;rain_draw[42][65] = 0;rain_draw[43][65] = 0;rain_draw[44][65] = 0;rain_draw[45][65] = 0;rain_draw[46][65] = 0;rain_draw[47][65] = 0;rain_draw[48][65] = 0;rain_draw[49][65] = 0;rain_draw[50][65] = 0;rain_draw[51][65] = 0;rain_draw[52][65] = 0;rain_draw[53][65] = 0;rain_draw[54][65] = 0;rain_draw[55][65] = 0;rain_draw[56][65] = 0;rain_draw[57][65] = 0;rain_draw[58][65] = 0;rain_draw[59][65] = 0;rain_draw[60][65] = 0;rain_draw[61][65] = 0;rain_draw[62][65] = 0;rain_draw[63][65] = 0;rain_draw[64][65] = 0;rain_draw[65][65] = 0;rain_draw[66][65] = 0;rain_draw[67][65] = 0;rain_draw[68][65] = 0;rain_draw[69][65] = 0;rain_draw[70][65] = 0;rain_draw[71][65] = 0;rain_draw[72][65] = 0;rain_draw[73][65] = 0;rain_draw[74][65] = 0;rain_draw[75][65] = 0;rain_draw[76][65] = 0;rain_draw[77][65] = 0;rain_draw[78][65] = 0;rain_draw[79][65] = 0;rain_draw[80][65] = 0;rain_draw[81][65] = 0;rain_draw[82][65] = 0;rain_draw[83][65] = 0;rain_draw[84][65] = 0;rain_draw[85][65] = 0;rain_draw[86][65] = 0;rain_draw[87][65] = 0;rain_draw[88][65] = 0;rain_draw[89][65] = 0;rain_draw[90][65] = 0;rain_draw[91][65] = 0;rain_draw[92][65] = 0;rain_draw[93][65] = 0;rain_draw[94][65] = 0;rain_draw[95][65] = 0;
        rain_draw[0][66] = 0;rain_draw[1][66] = 0;rain_draw[2][66] = 0;rain_draw[3][66] = 0;rain_draw[4][66] = 0;rain_draw[5][66] = 0;rain_draw[6][66] = 0;rain_draw[7][66] = 0;rain_draw[8][66] = 0;rain_draw[9][66] = 0;rain_draw[10][66] = 0;rain_draw[11][66] = 0;rain_draw[12][66] = 0;rain_draw[13][66] = 0;rain_draw[14][66] = 0;rain_draw[15][66] = 0;rain_draw[16][66] = 1;rain_draw[17][66] = 1;rain_draw[18][66] = 1;rain_draw[19][66] = 0;rain_draw[20][66] = 0;rain_draw[21][66] = 0;rain_draw[22][66] = 0;rain_draw[23][66] = 0;rain_draw[24][66] = 0;rain_draw[25][66] = 0;rain_draw[26][66] = 0;rain_draw[27][66] = 0;rain_draw[28][66] = 0;rain_draw[29][66] = 0;rain_draw[30][66] = 0;rain_draw[31][66] = 0;rain_draw[32][66] = 0;rain_draw[33][66] = 0;rain_draw[34][66] = 0;rain_draw[35][66] = 0;rain_draw[36][66] = 0;rain_draw[37][66] = 0;rain_draw[38][66] = 0;rain_draw[39][66] = 0;rain_draw[40][66] = 0;rain_draw[41][66] = 0;rain_draw[42][66] = 0;rain_draw[43][66] = 0;rain_draw[44][66] = 0;rain_draw[45][66] = 0;rain_draw[46][66] = 0;rain_draw[47][66] = 1;rain_draw[48][66] = 1;rain_draw[49][66] = 1;rain_draw[50][66] = 0;rain_draw[51][66] = 0;rain_draw[52][66] = 0;rain_draw[53][66] = 0;rain_draw[54][66] = 0;rain_draw[55][66] = 0;rain_draw[56][66] = 0;rain_draw[57][66] = 0;rain_draw[58][66] = 0;rain_draw[59][66] = 0;rain_draw[60][66] = 0;rain_draw[61][66] = 0;rain_draw[62][66] = 0;rain_draw[63][66] = 0;rain_draw[64][66] = 0;rain_draw[65][66] = 0;rain_draw[66][66] = 0;rain_draw[67][66] = 0;rain_draw[68][66] = 0;rain_draw[69][66] = 0;rain_draw[70][66] = 0;rain_draw[71][66] = 0;rain_draw[72][66] = 0;rain_draw[73][66] = 0;rain_draw[74][66] = 0;rain_draw[75][66] = 0;rain_draw[76][66] = 0;rain_draw[77][66] = 0;rain_draw[78][66] = 0;rain_draw[79][66] = 0;rain_draw[80][66] = 0;rain_draw[81][66] = 0;rain_draw[82][66] = 0;rain_draw[83][66] = 0;rain_draw[84][66] = 0;rain_draw[85][66] = 0;rain_draw[86][66] = 0;rain_draw[87][66] = 0;rain_draw[88][66] = 0;rain_draw[89][66] = 0;rain_draw[90][66] = 0;rain_draw[91][66] = 0;rain_draw[92][66] = 0;rain_draw[93][66] = 0;rain_draw[94][66] = 0;rain_draw[95][66] = 0;
        rain_draw[0][67] = 0;rain_draw[1][67] = 0;rain_draw[2][67] = 0;rain_draw[3][67] = 0;rain_draw[4][67] = 0;rain_draw[5][67] = 0;rain_draw[6][67] = 0;rain_draw[7][67] = 0;rain_draw[8][67] = 0;rain_draw[9][67] = 0;rain_draw[10][67] = 0;rain_draw[11][67] = 0;rain_draw[12][67] = 0;rain_draw[13][67] = 0;rain_draw[14][67] = 0;rain_draw[15][67] = 1;rain_draw[16][67] = 1;rain_draw[17][67] = 1;rain_draw[18][67] = 0;rain_draw[19][67] = 0;rain_draw[20][67] = 0;rain_draw[21][67] = 0;rain_draw[22][67] = 0;rain_draw[23][67] = 0;rain_draw[24][67] = 0;rain_draw[25][67] = 0;rain_draw[26][67] = 0;rain_draw[27][67] = 0;rain_draw[28][67] = 0;rain_draw[29][67] = 0;rain_draw[30][67] = 0;rain_draw[31][67] = 0;rain_draw[32][67] = 0;rain_draw[33][67] = 0;rain_draw[34][67] = 0;rain_draw[35][67] = 0;rain_draw[36][67] = 0;rain_draw[37][67] = 0;rain_draw[38][67] = 0;rain_draw[39][67] = 0;rain_draw[40][67] = 0;rain_draw[41][67] = 0;rain_draw[42][67] = 0;rain_draw[43][67] = 0;rain_draw[44][67] = 0;rain_draw[45][67] = 0;rain_draw[46][67] = 1;rain_draw[47][67] = 1;rain_draw[48][67] = 1;rain_draw[49][67] = 0;rain_draw[50][67] = 0;rain_draw[51][67] = 0;rain_draw[52][67] = 0;rain_draw[53][67] = 0;rain_draw[54][67] = 0;rain_draw[55][67] = 0;rain_draw[56][67] = 0;rain_draw[57][67] = 0;rain_draw[58][67] = 0;rain_draw[59][67] = 0;rain_draw[60][67] = 0;rain_draw[61][67] = 0;rain_draw[62][67] = 0;rain_draw[63][67] = 0;rain_draw[64][67] = 0;rain_draw[65][67] = 0;rain_draw[66][67] = 0;rain_draw[67][67] = 0;rain_draw[68][67] = 0;rain_draw[69][67] = 0;rain_draw[70][67] = 0;rain_draw[71][67] = 0;rain_draw[72][67] = 0;rain_draw[73][67] = 0;rain_draw[74][67] = 0;rain_draw[75][67] = 0;rain_draw[76][67] = 0;rain_draw[77][67] = 0;rain_draw[78][67] = 0;rain_draw[79][67] = 0;rain_draw[80][67] = 0;rain_draw[81][67] = 0;rain_draw[82][67] = 0;rain_draw[83][67] = 0;rain_draw[84][67] = 0;rain_draw[85][67] = 0;rain_draw[86][67] = 0;rain_draw[87][67] = 0;rain_draw[88][67] = 0;rain_draw[89][67] = 0;rain_draw[90][67] = 0;rain_draw[91][67] = 0;rain_draw[92][67] = 0;rain_draw[93][67] = 0;rain_draw[94][67] = 0;rain_draw[95][67] = 0;
        rain_draw[0][68] = 0;rain_draw[1][68] = 0;rain_draw[2][68] = 0;rain_draw[3][68] = 0;rain_draw[4][68] = 0;rain_draw[5][68] = 0;rain_draw[6][68] = 0;rain_draw[7][68] = 0;rain_draw[8][68] = 0;rain_draw[9][68] = 0;rain_draw[10][68] = 0;rain_draw[11][68] = 0;rain_draw[12][68] = 0;rain_draw[13][68] = 0;rain_draw[14][68] = 1;rain_draw[15][68] = 1;rain_draw[16][68] = 1;rain_draw[17][68] = 0;rain_draw[18][68] = 0;rain_draw[19][68] = 0;rain_draw[20][68] = 0;rain_draw[21][68] = 0;rain_draw[22][68] = 0;rain_draw[23][68] = 0;rain_draw[24][68] = 0;rain_draw[25][68] = 0;rain_draw[26][68] = 0;rain_draw[27][68] = 0;rain_draw[28][68] = 0;rain_draw[29][68] = 0;rain_draw[30][68] = 0;rain_draw[31][68] = 0;rain_draw[32][68] = 0;rain_draw[33][68] = 0;rain_draw[34][68] = 0;rain_draw[35][68] = 0;rain_draw[36][68] = 0;rain_draw[37][68] = 0;rain_draw[38][68] = 0;rain_draw[39][68] = 0;rain_draw[40][68] = 0;rain_draw[41][68] = 0;rain_draw[42][68] = 0;rain_draw[43][68] = 0;rain_draw[44][68] = 0;rain_draw[45][68] = 1;rain_draw[46][68] = 1;rain_draw[47][68] = 1;rain_draw[48][68] = 0;rain_draw[49][68] = 0;rain_draw[50][68] = 0;rain_draw[51][68] = 0;rain_draw[52][68] = 0;rain_draw[53][68] = 0;rain_draw[54][68] = 0;rain_draw[55][68] = 0;rain_draw[56][68] = 0;rain_draw[57][68] = 0;rain_draw[58][68] = 0;rain_draw[59][68] = 0;rain_draw[60][68] = 0;rain_draw[61][68] = 0;rain_draw[62][68] = 0;rain_draw[63][68] = 0;rain_draw[64][68] = 0;rain_draw[65][68] = 0;rain_draw[66][68] = 0;rain_draw[67][68] = 0;rain_draw[68][68] = 0;rain_draw[69][68] = 0;rain_draw[70][68] = 0;rain_draw[71][68] = 0;rain_draw[72][68] = 0;rain_draw[73][68] = 0;rain_draw[74][68] = 0;rain_draw[75][68] = 0;rain_draw[76][68] = 0;rain_draw[77][68] = 0;rain_draw[78][68] = 0;rain_draw[79][68] = 0;rain_draw[80][68] = 0;rain_draw[81][68] = 0;rain_draw[82][68] = 0;rain_draw[83][68] = 0;rain_draw[84][68] = 0;rain_draw[85][68] = 0;rain_draw[86][68] = 0;rain_draw[87][68] = 0;rain_draw[88][68] = 0;rain_draw[89][68] = 0;rain_draw[90][68] = 0;rain_draw[91][68] = 0;rain_draw[92][68] = 0;rain_draw[93][68] = 0;rain_draw[94][68] = 0;rain_draw[95][68] = 0;
        rain_draw[0][69] = 0;rain_draw[1][69] = 0;rain_draw[2][69] = 0;rain_draw[3][69] = 0;rain_draw[4][69] = 0;rain_draw[5][69] = 0;rain_draw[6][69] = 0;rain_draw[7][69] = 0;rain_draw[8][69] = 0;rain_draw[9][69] = 0;rain_draw[10][69] = 0;rain_draw[11][69] = 0;rain_draw[12][69] = 0;rain_draw[13][69] = 1;rain_draw[14][69] = 1;rain_draw[15][69] = 1;rain_draw[16][69] = 0;rain_draw[17][69] = 0;rain_draw[18][69] = 0;rain_draw[19][69] = 0;rain_draw[20][69] = 0;rain_draw[21][69] = 0;rain_draw[22][69] = 0;rain_draw[23][69] = 0;rain_draw[24][69] = 0;rain_draw[25][69] = 0;rain_draw[26][69] = 0;rain_draw[27][69] = 0;rain_draw[28][69] = 0;rain_draw[29][69] = 0;rain_draw[30][69] = 0;rain_draw[31][69] = 0;rain_draw[32][69] = 0;rain_draw[33][69] = 0;rain_draw[34][69] = 0;rain_draw[35][69] = 0;rain_draw[36][69] = 0;rain_draw[37][69] = 0;rain_draw[38][69] = 0;rain_draw[39][69] = 0;rain_draw[40][69] = 0;rain_draw[41][69] = 0;rain_draw[42][69] = 0;rain_draw[43][69] = 0;rain_draw[44][69] = 1;rain_draw[45][69] = 1;rain_draw[46][69] = 1;rain_draw[47][69] = 0;rain_draw[48][69] = 0;rain_draw[49][69] = 0;rain_draw[50][69] = 0;rain_draw[51][69] = 0;rain_draw[52][69] = 0;rain_draw[53][69] = 0;rain_draw[54][69] = 0;rain_draw[55][69] = 0;rain_draw[56][69] = 0;rain_draw[57][69] = 0;rain_draw[58][69] = 0;rain_draw[59][69] = 0;rain_draw[60][69] = 0;rain_draw[61][69] = 0;rain_draw[62][69] = 0;rain_draw[63][69] = 0;rain_draw[64][69] = 0;rain_draw[65][69] = 0;rain_draw[66][69] = 0;rain_draw[67][69] = 0;rain_draw[68][69] = 0;rain_draw[69][69] = 0;rain_draw[70][69] = 0;rain_draw[71][69] = 0;rain_draw[72][69] = 0;rain_draw[73][69] = 0;rain_draw[74][69] = 0;rain_draw[75][69] = 0;rain_draw[76][69] = 0;rain_draw[77][69] = 0;rain_draw[78][69] = 0;rain_draw[79][69] = 0;rain_draw[80][69] = 0;rain_draw[81][69] = 0;rain_draw[82][69] = 0;rain_draw[83][69] = 0;rain_draw[84][69] = 0;rain_draw[85][69] = 0;rain_draw[86][69] = 0;rain_draw[87][69] = 0;rain_draw[88][69] = 0;rain_draw[89][69] = 0;rain_draw[90][69] = 0;rain_draw[91][69] = 0;rain_draw[92][69] = 0;rain_draw[93][69] = 0;rain_draw[94][69] = 0;rain_draw[95][69] = 0;
        rain_draw[0][70] = 0;rain_draw[1][70] = 0;rain_draw[2][70] = 0;rain_draw[3][70] = 0;rain_draw[4][70] = 0;rain_draw[5][70] = 0;rain_draw[6][70] = 0;rain_draw[7][70] = 0;rain_draw[8][70] = 0;rain_draw[9][70] = 0;rain_draw[10][70] = 0;rain_draw[11][70] = 0;rain_draw[12][70] = 1;rain_draw[13][70] = 1;rain_draw[14][70] = 1;rain_draw[15][70] = 0;rain_draw[16][70] = 0;rain_draw[17][70] = 0;rain_draw[18][70] = 0;rain_draw[19][70] = 0;rain_draw[20][70] = 0;rain_draw[21][70] = 0;rain_draw[22][70] = 0;rain_draw[23][70] = 0;rain_draw[24][70] = 0;rain_draw[25][70] = 0;rain_draw[26][70] = 0;rain_draw[27][70] = 0;rain_draw[28][70] = 0;rain_draw[29][70] = 0;rain_draw[30][70] = 0;rain_draw[31][70] = 0;rain_draw[32][70] = 0;rain_draw[33][70] = 0;rain_draw[34][70] = 0;rain_draw[35][70] = 0;rain_draw[36][70] = 0;rain_draw[37][70] = 0;rain_draw[38][70] = 0;rain_draw[39][70] = 0;rain_draw[40][70] = 0;rain_draw[41][70] = 0;rain_draw[42][70] = 0;rain_draw[43][70] = 1;rain_draw[44][70] = 1;rain_draw[45][70] = 1;rain_draw[46][70] = 0;rain_draw[47][70] = 0;rain_draw[48][70] = 0;rain_draw[49][70] = 0;rain_draw[50][70] = 0;rain_draw[51][70] = 0;rain_draw[52][70] = 0;rain_draw[53][70] = 0;rain_draw[54][70] = 0;rain_draw[55][70] = 0;rain_draw[56][70] = 0;rain_draw[57][70] = 0;rain_draw[58][70] = 0;rain_draw[59][70] = 0;rain_draw[60][70] = 0;rain_draw[61][70] = 0;rain_draw[62][70] = 0;rain_draw[63][70] = 0;rain_draw[64][70] = 0;rain_draw[65][70] = 0;rain_draw[66][70] = 0;rain_draw[67][70] = 0;rain_draw[68][70] = 0;rain_draw[69][70] = 0;rain_draw[70][70] = 0;rain_draw[71][70] = 0;rain_draw[72][70] = 0;rain_draw[73][70] = 0;rain_draw[74][70] = 0;rain_draw[75][70] = 0;rain_draw[76][70] = 0;rain_draw[77][70] = 0;rain_draw[78][70] = 0;rain_draw[79][70] = 0;rain_draw[80][70] = 0;rain_draw[81][70] = 0;rain_draw[82][70] = 0;rain_draw[83][70] = 0;rain_draw[84][70] = 0;rain_draw[85][70] = 0;rain_draw[86][70] = 0;rain_draw[87][70] = 0;rain_draw[88][70] = 0;rain_draw[89][70] = 0;rain_draw[90][70] = 0;rain_draw[91][70] = 0;rain_draw[92][70] = 0;rain_draw[93][70] = 0;rain_draw[94][70] = 0;rain_draw[95][70] = 0;
        rain_draw[0][71] = 0;rain_draw[1][71] = 0;rain_draw[2][71] = 0;rain_draw[3][71] = 0;rain_draw[4][71] = 0;rain_draw[5][71] = 0;rain_draw[6][71] = 0;rain_draw[7][71] = 0;rain_draw[8][71] = 0;rain_draw[9][71] = 0;rain_draw[10][71] = 0;rain_draw[11][71] = 1;rain_draw[12][71] = 1;rain_draw[13][71] = 1;rain_draw[14][71] = 0;rain_draw[15][71] = 0;rain_draw[16][71] = 0;rain_draw[17][71] = 0;rain_draw[18][71] = 0;rain_draw[19][71] = 0;rain_draw[20][71] = 0;rain_draw[21][71] = 0;rain_draw[22][71] = 0;rain_draw[23][71] = 0;rain_draw[24][71] = 0;rain_draw[25][71] = 0;rain_draw[26][71] = 0;rain_draw[27][71] = 0;rain_draw[28][71] = 0;rain_draw[29][71] = 0;rain_draw[30][71] = 0;rain_draw[31][71] = 0;rain_draw[32][71] = 0;rain_draw[33][71] = 0;rain_draw[34][71] = 0;rain_draw[35][71] = 0;rain_draw[36][71] = 0;rain_draw[37][71] = 0;rain_draw[38][71] = 0;rain_draw[39][71] = 0;rain_draw[40][71] = 0;rain_draw[41][71] = 0;rain_draw[42][71] = 1;rain_draw[43][71] = 1;rain_draw[44][71] = 1;rain_draw[45][71] = 0;rain_draw[46][71] = 0;rain_draw[47][71] = 0;rain_draw[48][71] = 0;rain_draw[49][71] = 0;rain_draw[50][71] = 0;rain_draw[51][71] = 0;rain_draw[52][71] = 0;rain_draw[53][71] = 0;rain_draw[54][71] = 0;rain_draw[55][71] = 0;rain_draw[56][71] = 0;rain_draw[57][71] = 0;rain_draw[58][71] = 0;rain_draw[59][71] = 0;rain_draw[60][71] = 0;rain_draw[61][71] = 0;rain_draw[62][71] = 0;rain_draw[63][71] = 0;rain_draw[64][71] = 0;rain_draw[65][71] = 0;rain_draw[66][71] = 0;rain_draw[67][71] = 0;rain_draw[68][71] = 0;rain_draw[69][71] = 0;rain_draw[70][71] = 0;rain_draw[71][71] = 0;rain_draw[72][71] = 0;rain_draw[73][71] = 0;rain_draw[74][71] = 0;rain_draw[75][71] = 0;rain_draw[76][71] = 0;rain_draw[77][71] = 0;rain_draw[78][71] = 0;rain_draw[79][71] = 0;rain_draw[80][71] = 0;rain_draw[81][71] = 0;rain_draw[82][71] = 0;rain_draw[83][71] = 0;rain_draw[84][71] = 0;rain_draw[85][71] = 0;rain_draw[86][71] = 0;rain_draw[87][71] = 0;rain_draw[88][71] = 0;rain_draw[89][71] = 0;rain_draw[90][71] = 0;rain_draw[91][71] = 0;rain_draw[92][71] = 0;rain_draw[93][71] = 0;rain_draw[94][71] = 0;rain_draw[95][71] = 0;
        rain_draw[0][72] = 0;rain_draw[1][72] = 0;rain_draw[2][72] = 0;rain_draw[3][72] = 0;rain_draw[4][72] = 0;rain_draw[5][72] = 0;rain_draw[6][72] = 0;rain_draw[7][72] = 0;rain_draw[8][72] = 0;rain_draw[9][72] = 0;rain_draw[10][72] = 1;rain_draw[11][72] = 1;rain_draw[12][72] = 1;rain_draw[13][72] = 0;rain_draw[14][72] = 0;rain_draw[15][72] = 0;rain_draw[16][72] = 0;rain_draw[17][72] = 0;rain_draw[18][72] = 0;rain_draw[19][72] = 0;rain_draw[20][72] = 0;rain_draw[21][72] = 0;rain_draw[22][72] = 0;rain_draw[23][72] = 0;rain_draw[24][72] = 0;rain_draw[25][72] = 0;rain_draw[26][72] = 0;rain_draw[27][72] = 0;rain_draw[28][72] = 0;rain_draw[29][72] = 0;rain_draw[30][72] = 0;rain_draw[31][72] = 0;rain_draw[32][72] = 0;rain_draw[33][72] = 0;rain_draw[34][72] = 0;rain_draw[35][72] = 0;rain_draw[36][72] = 0;rain_draw[37][72] = 0;rain_draw[38][72] = 0;rain_draw[39][72] = 0;rain_draw[40][72] = 0;rain_draw[41][72] = 1;rain_draw[42][72] = 1;rain_draw[43][72] = 1;rain_draw[44][72] = 0;rain_draw[45][72] = 0;rain_draw[46][72] = 0;rain_draw[47][72] = 0;rain_draw[48][72] = 0;rain_draw[49][72] = 0;rain_draw[50][72] = 0;rain_draw[51][72] = 0;rain_draw[52][72] = 0;rain_draw[53][72] = 0;rain_draw[54][72] = 0;rain_draw[55][72] = 0;rain_draw[56][72] = 0;rain_draw[57][72] = 0;rain_draw[58][72] = 0;rain_draw[59][72] = 0;rain_draw[60][72] = 0;rain_draw[61][72] = 0;rain_draw[62][72] = 0;rain_draw[63][72] = 0;rain_draw[64][72] = 0;rain_draw[65][72] = 0;rain_draw[66][72] = 0;rain_draw[67][72] = 0;rain_draw[68][72] = 0;rain_draw[69][72] = 0;rain_draw[70][72] = 0;rain_draw[71][72] = 0;rain_draw[72][72] = 0;rain_draw[73][72] = 0;rain_draw[74][72] = 0;rain_draw[75][72] = 0;rain_draw[76][72] = 0;rain_draw[77][72] = 0;rain_draw[78][72] = 0;rain_draw[79][72] = 0;rain_draw[80][72] = 0;rain_draw[81][72] = 0;rain_draw[82][72] = 0;rain_draw[83][72] = 0;rain_draw[84][72] = 0;rain_draw[85][72] = 0;rain_draw[86][72] = 0;rain_draw[87][72] = 0;rain_draw[88][72] = 0;rain_draw[89][72] = 0;rain_draw[90][72] = 0;rain_draw[91][72] = 0;rain_draw[92][72] = 0;rain_draw[93][72] = 0;rain_draw[94][72] = 0;rain_draw[95][72] = 0;
        rain_draw[0][73] = 0;rain_draw[1][73] = 0;rain_draw[2][73] = 0;rain_draw[3][73] = 0;rain_draw[4][73] = 0;rain_draw[5][73] = 0;rain_draw[6][73] = 0;rain_draw[7][73] = 0;rain_draw[8][73] = 0;rain_draw[9][73] = 0;rain_draw[10][73] = 0;rain_draw[11][73] = 0;rain_draw[12][73] = 0;rain_draw[13][73] = 0;rain_draw[14][73] = 0;rain_draw[15][73] = 0;rain_draw[16][73] = 0;rain_draw[17][73] = 0;rain_draw[18][73] = 0;rain_draw[19][73] = 0;rain_draw[20][73] = 0;rain_draw[21][73] = 0;rain_draw[22][73] = 0;rain_draw[23][73] = 0;rain_draw[24][73] = 0;rain_draw[25][73] = 0;rain_draw[26][73] = 0;rain_draw[27][73] = 0;rain_draw[28][73] = 0;rain_draw[29][73] = 0;rain_draw[30][73] = 0;rain_draw[31][73] = 0;rain_draw[32][73] = 0;rain_draw[33][73] = 0;rain_draw[34][73] = 0;rain_draw[35][73] = 0;rain_draw[36][73] = 0;rain_draw[37][73] = 0;rain_draw[38][73] = 0;rain_draw[39][73] = 0;rain_draw[40][73] = 0;rain_draw[41][73] = 0;rain_draw[42][73] = 0;rain_draw[43][73] = 0;rain_draw[44][73] = 0;rain_draw[45][73] = 0;rain_draw[46][73] = 0;rain_draw[47][73] = 0;rain_draw[48][73] = 0;rain_draw[49][73] = 0;rain_draw[50][73] = 0;rain_draw[51][73] = 0;rain_draw[52][73] = 0;rain_draw[53][73] = 0;rain_draw[54][73] = 0;rain_draw[55][73] = 0;rain_draw[56][73] = 0;rain_draw[57][73] = 0;rain_draw[58][73] = 0;rain_draw[59][73] = 0;rain_draw[60][73] = 0;rain_draw[61][73] = 0;rain_draw[62][73] = 0;rain_draw[63][73] = 0;rain_draw[64][73] = 0;rain_draw[65][73] = 0;rain_draw[66][73] = 0;rain_draw[67][73] = 0;rain_draw[68][73] = 0;rain_draw[69][73] = 0;rain_draw[70][73] = 0;rain_draw[71][73] = 0;rain_draw[72][73] = 0;rain_draw[73][73] = 0;rain_draw[74][73] = 0;rain_draw[75][73] = 0;rain_draw[76][73] = 0;rain_draw[77][73] = 0;rain_draw[78][73] = 0;rain_draw[79][73] = 0;rain_draw[80][73] = 0;rain_draw[81][73] = 0;rain_draw[82][73] = 0;rain_draw[83][73] = 0;rain_draw[84][73] = 0;rain_draw[85][73] = 0;rain_draw[86][73] = 0;rain_draw[87][73] = 0;rain_draw[88][73] = 0;rain_draw[89][73] = 0;rain_draw[90][73] = 0;rain_draw[91][73] = 0;rain_draw[92][73] = 0;rain_draw[93][73] = 0;rain_draw[94][73] = 0;rain_draw[95][73] = 0;
        rain_draw[0][74] = 0;rain_draw[1][74] = 0;rain_draw[2][74] = 0;rain_draw[3][74] = 0;rain_draw[4][74] = 0;rain_draw[5][74] = 0;rain_draw[6][74] = 0;rain_draw[7][74] = 0;rain_draw[8][74] = 0;rain_draw[9][74] = 0;rain_draw[10][74] = 0;rain_draw[11][74] = 0;rain_draw[12][74] = 0;rain_draw[13][74] = 0;rain_draw[14][74] = 0;rain_draw[15][74] = 0;rain_draw[16][74] = 0;rain_draw[17][74] = 0;rain_draw[18][74] = 0;rain_draw[19][74] = 0;rain_draw[20][74] = 0;rain_draw[21][74] = 0;rain_draw[22][74] = 0;rain_draw[23][74] = 0;rain_draw[24][74] = 0;rain_draw[25][74] = 0;rain_draw[26][74] = 0;rain_draw[27][74] = 0;rain_draw[28][74] = 0;rain_draw[29][74] = 0;rain_draw[30][74] = 0;rain_draw[31][74] = 0;rain_draw[32][74] = 0;rain_draw[33][74] = 0;rain_draw[34][74] = 0;rain_draw[35][74] = 0;rain_draw[36][74] = 0;rain_draw[37][74] = 0;rain_draw[38][74] = 0;rain_draw[39][74] = 0;rain_draw[40][74] = 0;rain_draw[41][74] = 0;rain_draw[42][74] = 0;rain_draw[43][74] = 0;rain_draw[44][74] = 0;rain_draw[45][74] = 0;rain_draw[46][74] = 0;rain_draw[47][74] = 0;rain_draw[48][74] = 0;rain_draw[49][74] = 0;rain_draw[50][74] = 0;rain_draw[51][74] = 0;rain_draw[52][74] = 0;rain_draw[53][74] = 0;rain_draw[54][74] = 0;rain_draw[55][74] = 0;rain_draw[56][74] = 0;rain_draw[57][74] = 0;rain_draw[58][74] = 0;rain_draw[59][74] = 0;rain_draw[60][74] = 0;rain_draw[61][74] = 0;rain_draw[62][74] = 0;rain_draw[63][74] = 0;rain_draw[64][74] = 0;rain_draw[65][74] = 0;rain_draw[66][74] = 0;rain_draw[67][74] = 0;rain_draw[68][74] = 0;rain_draw[69][74] = 0;rain_draw[70][74] = 0;rain_draw[71][74] = 0;rain_draw[72][74] = 0;rain_draw[73][74] = 0;rain_draw[74][74] = 0;rain_draw[75][74] = 0;rain_draw[76][74] = 0;rain_draw[77][74] = 0;rain_draw[78][74] = 0;rain_draw[79][74] = 0;rain_draw[80][74] = 0;rain_draw[81][74] = 0;rain_draw[82][74] = 0;rain_draw[83][74] = 0;rain_draw[84][74] = 0;rain_draw[85][74] = 0;rain_draw[86][74] = 0;rain_draw[87][74] = 0;rain_draw[88][74] = 0;rain_draw[89][74] = 0;rain_draw[90][74] = 0;rain_draw[91][74] = 0;rain_draw[92][74] = 0;rain_draw[93][74] = 0;rain_draw[94][74] = 0;rain_draw[95][74] = 0;
        rain_draw[0][75] = 0;rain_draw[1][75] = 0;rain_draw[2][75] = 0;rain_draw[3][75] = 0;rain_draw[4][75] = 0;rain_draw[5][75] = 0;rain_draw[6][75] = 0;rain_draw[7][75] = 0;rain_draw[8][75] = 0;rain_draw[9][75] = 0;rain_draw[10][75] = 0;rain_draw[11][75] = 0;rain_draw[12][75] = 0;rain_draw[13][75] = 0;rain_draw[14][75] = 0;rain_draw[15][75] = 0;rain_draw[16][75] = 0;rain_draw[17][75] = 0;rain_draw[18][75] = 0;rain_draw[19][75] = 0;rain_draw[20][75] = 0;rain_draw[21][75] = 0;rain_draw[22][75] = 0;rain_draw[23][75] = 0;rain_draw[24][75] = 0;rain_draw[25][75] = 0;rain_draw[26][75] = 0;rain_draw[27][75] = 0;rain_draw[28][75] = 0;rain_draw[29][75] = 0;rain_draw[30][75] = 0;rain_draw[31][75] = 0;rain_draw[32][75] = 0;rain_draw[33][75] = 0;rain_draw[34][75] = 0;rain_draw[35][75] = 0;rain_draw[36][75] = 0;rain_draw[37][75] = 0;rain_draw[38][75] = 0;rain_draw[39][75] = 0;rain_draw[40][75] = 0;rain_draw[41][75] = 0;rain_draw[42][75] = 0;rain_draw[43][75] = 0;rain_draw[44][75] = 0;rain_draw[45][75] = 0;rain_draw[46][75] = 0;rain_draw[47][75] = 0;rain_draw[48][75] = 0;rain_draw[49][75] = 0;rain_draw[50][75] = 0;rain_draw[51][75] = 0;rain_draw[52][75] = 0;rain_draw[53][75] = 0;rain_draw[54][75] = 0;rain_draw[55][75] = 0;rain_draw[56][75] = 0;rain_draw[57][75] = 0;rain_draw[58][75] = 0;rain_draw[59][75] = 0;rain_draw[60][75] = 0;rain_draw[61][75] = 0;rain_draw[62][75] = 0;rain_draw[63][75] = 0;rain_draw[64][75] = 0;rain_draw[65][75] = 0;rain_draw[66][75] = 0;rain_draw[67][75] = 0;rain_draw[68][75] = 1;rain_draw[69][75] = 1;rain_draw[70][75] = 1;rain_draw[71][75] = 0;rain_draw[72][75] = 0;rain_draw[73][75] = 0;rain_draw[74][75] = 0;rain_draw[75][75] = 0;rain_draw[76][75] = 0;rain_draw[77][75] = 0;rain_draw[78][75] = 0;rain_draw[79][75] = 0;rain_draw[80][75] = 0;rain_draw[81][75] = 0;rain_draw[82][75] = 0;rain_draw[83][75] = 0;rain_draw[84][75] = 0;rain_draw[85][75] = 0;rain_draw[86][75] = 0;rain_draw[87][75] = 0;rain_draw[88][75] = 0;rain_draw[89][75] = 0;rain_draw[90][75] = 0;rain_draw[91][75] = 0;rain_draw[92][75] = 0;rain_draw[93][75] = 0;rain_draw[94][75] = 0;rain_draw[95][75] = 0;
        rain_draw[0][76] = 0;rain_draw[1][76] = 0;rain_draw[2][76] = 0;rain_draw[3][76] = 0;rain_draw[4][76] = 0;rain_draw[5][76] = 0;rain_draw[6][76] = 0;rain_draw[7][76] = 0;rain_draw[8][76] = 0;rain_draw[9][76] = 0;rain_draw[10][76] = 0;rain_draw[11][76] = 0;rain_draw[12][76] = 0;rain_draw[13][76] = 0;rain_draw[14][76] = 0;rain_draw[15][76] = 0;rain_draw[16][76] = 0;rain_draw[17][76] = 0;rain_draw[18][76] = 0;rain_draw[19][76] = 0;rain_draw[20][76] = 0;rain_draw[21][76] = 0;rain_draw[22][76] = 0;rain_draw[23][76] = 0;rain_draw[24][76] = 0;rain_draw[25][76] = 0;rain_draw[26][76] = 0;rain_draw[27][76] = 0;rain_draw[28][76] = 0;rain_draw[29][76] = 0;rain_draw[30][76] = 0;rain_draw[31][76] = 0;rain_draw[32][76] = 0;rain_draw[33][76] = 0;rain_draw[34][76] = 0;rain_draw[35][76] = 0;rain_draw[36][76] = 0;rain_draw[37][76] = 0;rain_draw[38][76] = 0;rain_draw[39][76] = 0;rain_draw[40][76] = 0;rain_draw[41][76] = 0;rain_draw[42][76] = 0;rain_draw[43][76] = 0;rain_draw[44][76] = 0;rain_draw[45][76] = 0;rain_draw[46][76] = 0;rain_draw[47][76] = 0;rain_draw[48][76] = 0;rain_draw[49][76] = 0;rain_draw[50][76] = 0;rain_draw[51][76] = 0;rain_draw[52][76] = 0;rain_draw[53][76] = 0;rain_draw[54][76] = 0;rain_draw[55][76] = 0;rain_draw[56][76] = 0;rain_draw[57][76] = 0;rain_draw[58][76] = 0;rain_draw[59][76] = 0;rain_draw[60][76] = 0;rain_draw[61][76] = 0;rain_draw[62][76] = 0;rain_draw[63][76] = 0;rain_draw[64][76] = 0;rain_draw[65][76] = 0;rain_draw[66][76] = 0;rain_draw[67][76] = 1;rain_draw[68][76] = 1;rain_draw[69][76] = 1;rain_draw[70][76] = 0;rain_draw[71][76] = 0;rain_draw[72][76] = 0;rain_draw[73][76] = 0;rain_draw[74][76] = 0;rain_draw[75][76] = 0;rain_draw[76][76] = 0;rain_draw[77][76] = 0;rain_draw[78][76] = 0;rain_draw[79][76] = 0;rain_draw[80][76] = 0;rain_draw[81][76] = 0;rain_draw[82][76] = 0;rain_draw[83][76] = 0;rain_draw[84][76] = 0;rain_draw[85][76] = 0;rain_draw[86][76] = 0;rain_draw[87][76] = 0;rain_draw[88][76] = 0;rain_draw[89][76] = 0;rain_draw[90][76] = 0;rain_draw[91][76] = 0;rain_draw[92][76] = 0;rain_draw[93][76] = 0;rain_draw[94][76] = 0;rain_draw[95][76] = 0;
        rain_draw[0][77] = 0;rain_draw[1][77] = 0;rain_draw[2][77] = 0;rain_draw[3][77] = 0;rain_draw[4][77] = 0;rain_draw[5][77] = 0;rain_draw[6][77] = 0;rain_draw[7][77] = 0;rain_draw[8][77] = 0;rain_draw[9][77] = 0;rain_draw[10][77] = 0;rain_draw[11][77] = 0;rain_draw[12][77] = 0;rain_draw[13][77] = 0;rain_draw[14][77] = 0;rain_draw[15][77] = 0;rain_draw[16][77] = 0;rain_draw[17][77] = 0;rain_draw[18][77] = 0;rain_draw[19][77] = 0;rain_draw[20][77] = 0;rain_draw[21][77] = 0;rain_draw[22][77] = 0;rain_draw[23][77] = 0;rain_draw[24][77] = 0;rain_draw[25][77] = 0;rain_draw[26][77] = 0;rain_draw[27][77] = 0;rain_draw[28][77] = 0;rain_draw[29][77] = 0;rain_draw[30][77] = 0;rain_draw[31][77] = 0;rain_draw[32][77] = 0;rain_draw[33][77] = 0;rain_draw[34][77] = 0;rain_draw[35][77] = 0;rain_draw[36][77] = 0;rain_draw[37][77] = 0;rain_draw[38][77] = 0;rain_draw[39][77] = 0;rain_draw[40][77] = 0;rain_draw[41][77] = 0;rain_draw[42][77] = 0;rain_draw[43][77] = 0;rain_draw[44][77] = 0;rain_draw[45][77] = 0;rain_draw[46][77] = 0;rain_draw[47][77] = 0;rain_draw[48][77] = 0;rain_draw[49][77] = 0;rain_draw[50][77] = 0;rain_draw[51][77] = 0;rain_draw[52][77] = 0;rain_draw[53][77] = 0;rain_draw[54][77] = 0;rain_draw[55][77] = 0;rain_draw[56][77] = 0;rain_draw[57][77] = 0;rain_draw[58][77] = 0;rain_draw[59][77] = 0;rain_draw[60][77] = 0;rain_draw[61][77] = 0;rain_draw[62][77] = 0;rain_draw[63][77] = 0;rain_draw[64][77] = 0;rain_draw[65][77] = 0;rain_draw[66][77] = 1;rain_draw[67][77] = 1;rain_draw[68][77] = 1;rain_draw[69][77] = 0;rain_draw[70][77] = 0;rain_draw[71][77] = 0;rain_draw[72][77] = 0;rain_draw[73][77] = 0;rain_draw[74][77] = 0;rain_draw[75][77] = 0;rain_draw[76][77] = 0;rain_draw[77][77] = 0;rain_draw[78][77] = 0;rain_draw[79][77] = 0;rain_draw[80][77] = 0;rain_draw[81][77] = 0;rain_draw[82][77] = 0;rain_draw[83][77] = 0;rain_draw[84][77] = 0;rain_draw[85][77] = 0;rain_draw[86][77] = 0;rain_draw[87][77] = 0;rain_draw[88][77] = 0;rain_draw[89][77] = 0;rain_draw[90][77] = 0;rain_draw[91][77] = 0;rain_draw[92][77] = 0;rain_draw[93][77] = 0;rain_draw[94][77] = 0;rain_draw[95][77] = 0;
        rain_draw[0][78] = 0;rain_draw[1][78] = 0;rain_draw[2][78] = 0;rain_draw[3][78] = 0;rain_draw[4][78] = 0;rain_draw[5][78] = 0;rain_draw[6][78] = 0;rain_draw[7][78] = 0;rain_draw[8][78] = 0;rain_draw[9][78] = 0;rain_draw[10][78] = 0;rain_draw[11][78] = 0;rain_draw[12][78] = 0;rain_draw[13][78] = 0;rain_draw[14][78] = 0;rain_draw[15][78] = 0;rain_draw[16][78] = 0;rain_draw[17][78] = 0;rain_draw[18][78] = 0;rain_draw[19][78] = 0;rain_draw[20][78] = 0;rain_draw[21][78] = 0;rain_draw[22][78] = 0;rain_draw[23][78] = 0;rain_draw[24][78] = 0;rain_draw[25][78] = 0;rain_draw[26][78] = 0;rain_draw[27][78] = 0;rain_draw[28][78] = 0;rain_draw[29][78] = 0;rain_draw[30][78] = 0;rain_draw[31][78] = 0;rain_draw[32][78] = 0;rain_draw[33][78] = 0;rain_draw[34][78] = 0;rain_draw[35][78] = 0;rain_draw[36][78] = 0;rain_draw[37][78] = 0;rain_draw[38][78] = 0;rain_draw[39][78] = 0;rain_draw[40][78] = 0;rain_draw[41][78] = 0;rain_draw[42][78] = 0;rain_draw[43][78] = 0;rain_draw[44][78] = 0;rain_draw[45][78] = 0;rain_draw[46][78] = 0;rain_draw[47][78] = 0;rain_draw[48][78] = 0;rain_draw[49][78] = 0;rain_draw[50][78] = 0;rain_draw[51][78] = 0;rain_draw[52][78] = 0;rain_draw[53][78] = 0;rain_draw[54][78] = 0;rain_draw[55][78] = 0;rain_draw[56][78] = 0;rain_draw[57][78] = 0;rain_draw[58][78] = 0;rain_draw[59][78] = 0;rain_draw[60][78] = 0;rain_draw[61][78] = 0;rain_draw[62][78] = 0;rain_draw[63][78] = 0;rain_draw[64][78] = 0;rain_draw[65][78] = 1;rain_draw[66][78] = 1;rain_draw[67][78] = 1;rain_draw[68][78] = 0;rain_draw[69][78] = 0;rain_draw[70][78] = 0;rain_draw[71][78] = 0;rain_draw[72][78] = 0;rain_draw[73][78] = 0;rain_draw[74][78] = 0;rain_draw[75][78] = 0;rain_draw[76][78] = 0;rain_draw[77][78] = 0;rain_draw[78][78] = 0;rain_draw[79][78] = 0;rain_draw[80][78] = 0;rain_draw[81][78] = 0;rain_draw[82][78] = 0;rain_draw[83][78] = 0;rain_draw[84][78] = 0;rain_draw[85][78] = 0;rain_draw[86][78] = 0;rain_draw[87][78] = 0;rain_draw[88][78] = 0;rain_draw[89][78] = 0;rain_draw[90][78] = 0;rain_draw[91][78] = 0;rain_draw[92][78] = 0;rain_draw[93][78] = 0;rain_draw[94][78] = 0;rain_draw[95][78] = 0;
        rain_draw[0][79] = 0;rain_draw[1][79] = 0;rain_draw[2][79] = 0;rain_draw[3][79] = 0;rain_draw[4][79] = 0;rain_draw[5][79] = 0;rain_draw[6][79] = 0;rain_draw[7][79] = 0;rain_draw[8][79] = 0;rain_draw[9][79] = 0;rain_draw[10][79] = 0;rain_draw[11][79] = 0;rain_draw[12][79] = 0;rain_draw[13][79] = 0;rain_draw[14][79] = 0;rain_draw[15][79] = 0;rain_draw[16][79] = 0;rain_draw[17][79] = 0;rain_draw[18][79] = 0;rain_draw[19][79] = 0;rain_draw[20][79] = 0;rain_draw[21][79] = 0;rain_draw[22][79] = 0;rain_draw[23][79] = 0;rain_draw[24][79] = 0;rain_draw[25][79] = 0;rain_draw[26][79] = 0;rain_draw[27][79] = 0;rain_draw[28][79] = 0;rain_draw[29][79] = 0;rain_draw[30][79] = 0;rain_draw[31][79] = 0;rain_draw[32][79] = 0;rain_draw[33][79] = 0;rain_draw[34][79] = 0;rain_draw[35][79] = 0;rain_draw[36][79] = 0;rain_draw[37][79] = 0;rain_draw[38][79] = 0;rain_draw[39][79] = 0;rain_draw[40][79] = 0;rain_draw[41][79] = 0;rain_draw[42][79] = 0;rain_draw[43][79] = 0;rain_draw[44][79] = 0;rain_draw[45][79] = 0;rain_draw[46][79] = 0;rain_draw[47][79] = 0;rain_draw[48][79] = 0;rain_draw[49][79] = 0;rain_draw[50][79] = 0;rain_draw[51][79] = 0;rain_draw[52][79] = 0;rain_draw[53][79] = 0;rain_draw[54][79] = 0;rain_draw[55][79] = 0;rain_draw[56][79] = 0;rain_draw[57][79] = 0;rain_draw[58][79] = 0;rain_draw[59][79] = 0;rain_draw[60][79] = 0;rain_draw[61][79] = 0;rain_draw[62][79] = 0;rain_draw[63][79] = 0;rain_draw[64][79] = 1;rain_draw[65][79] = 1;rain_draw[66][79] = 1;rain_draw[67][79] = 0;rain_draw[68][79] = 0;rain_draw[69][79] = 0;rain_draw[70][79] = 0;rain_draw[71][79] = 0;rain_draw[72][79] = 0;rain_draw[73][79] = 0;rain_draw[74][79] = 0;rain_draw[75][79] = 0;rain_draw[76][79] = 0;rain_draw[77][79] = 0;rain_draw[78][79] = 0;rain_draw[79][79] = 0;rain_draw[80][79] = 0;rain_draw[81][79] = 0;rain_draw[82][79] = 0;rain_draw[83][79] = 0;rain_draw[84][79] = 0;rain_draw[85][79] = 0;rain_draw[86][79] = 0;rain_draw[87][79] = 0;rain_draw[88][79] = 0;rain_draw[89][79] = 0;rain_draw[90][79] = 0;rain_draw[91][79] = 0;rain_draw[92][79] = 0;rain_draw[93][79] = 0;rain_draw[94][79] = 0;rain_draw[95][79] = 0;
        rain_draw[0][80] = 0;rain_draw[1][80] = 0;rain_draw[2][80] = 0;rain_draw[3][80] = 0;rain_draw[4][80] = 0;rain_draw[5][80] = 0;rain_draw[6][80] = 0;rain_draw[7][80] = 0;rain_draw[8][80] = 0;rain_draw[9][80] = 0;rain_draw[10][80] = 0;rain_draw[11][80] = 0;rain_draw[12][80] = 0;rain_draw[13][80] = 0;rain_draw[14][80] = 0;rain_draw[15][80] = 0;rain_draw[16][80] = 0;rain_draw[17][80] = 0;rain_draw[18][80] = 0;rain_draw[19][80] = 0;rain_draw[20][80] = 0;rain_draw[21][80] = 0;rain_draw[22][80] = 0;rain_draw[23][80] = 0;rain_draw[24][80] = 0;rain_draw[25][80] = 0;rain_draw[26][80] = 0;rain_draw[27][80] = 0;rain_draw[28][80] = 0;rain_draw[29][80] = 1;rain_draw[30][80] = 1;rain_draw[31][80] = 1;rain_draw[32][80] = 0;rain_draw[33][80] = 0;rain_draw[34][80] = 0;rain_draw[35][80] = 0;rain_draw[36][80] = 0;rain_draw[37][80] = 0;rain_draw[38][80] = 0;rain_draw[39][80] = 0;rain_draw[40][80] = 0;rain_draw[41][80] = 0;rain_draw[42][80] = 0;rain_draw[43][80] = 0;rain_draw[44][80] = 0;rain_draw[45][80] = 0;rain_draw[46][80] = 0;rain_draw[47][80] = 0;rain_draw[48][80] = 0;rain_draw[49][80] = 0;rain_draw[50][80] = 0;rain_draw[51][80] = 0;rain_draw[52][80] = 0;rain_draw[53][80] = 0;rain_draw[54][80] = 0;rain_draw[55][80] = 0;rain_draw[56][80] = 0;rain_draw[57][80] = 0;rain_draw[58][80] = 0;rain_draw[59][80] = 0;rain_draw[60][80] = 0;rain_draw[61][80] = 0;rain_draw[62][80] = 0;rain_draw[63][80] = 1;rain_draw[64][80] = 1;rain_draw[65][80] = 1;rain_draw[66][80] = 0;rain_draw[67][80] = 0;rain_draw[68][80] = 0;rain_draw[69][80] = 0;rain_draw[70][80] = 0;rain_draw[71][80] = 0;rain_draw[72][80] = 0;rain_draw[73][80] = 0;rain_draw[74][80] = 0;rain_draw[75][80] = 0;rain_draw[76][80] = 0;rain_draw[77][80] = 0;rain_draw[78][80] = 0;rain_draw[79][80] = 0;rain_draw[80][80] = 0;rain_draw[81][80] = 0;rain_draw[82][80] = 0;rain_draw[83][80] = 0;rain_draw[84][80] = 0;rain_draw[85][80] = 0;rain_draw[86][80] = 0;rain_draw[87][80] = 0;rain_draw[88][80] = 0;rain_draw[89][80] = 0;rain_draw[90][80] = 0;rain_draw[91][80] = 0;rain_draw[92][80] = 0;rain_draw[93][80] = 0;rain_draw[94][80] = 0;rain_draw[95][80] = 0;
        rain_draw[0][81] = 0;rain_draw[1][81] = 0;rain_draw[2][81] = 0;rain_draw[3][81] = 0;rain_draw[4][81] = 0;rain_draw[5][81] = 0;rain_draw[6][81] = 0;rain_draw[7][81] = 0;rain_draw[8][81] = 0;rain_draw[9][81] = 0;rain_draw[10][81] = 0;rain_draw[11][81] = 0;rain_draw[12][81] = 0;rain_draw[13][81] = 0;rain_draw[14][81] = 0;rain_draw[15][81] = 0;rain_draw[16][81] = 0;rain_draw[17][81] = 0;rain_draw[18][81] = 0;rain_draw[19][81] = 0;rain_draw[20][81] = 0;rain_draw[21][81] = 0;rain_draw[22][81] = 0;rain_draw[23][81] = 0;rain_draw[24][81] = 0;rain_draw[25][81] = 0;rain_draw[26][81] = 0;rain_draw[27][81] = 0;rain_draw[28][81] = 1;rain_draw[29][81] = 1;rain_draw[30][81] = 1;rain_draw[31][81] = 0;rain_draw[32][81] = 0;rain_draw[33][81] = 0;rain_draw[34][81] = 0;rain_draw[35][81] = 0;rain_draw[36][81] = 0;rain_draw[37][81] = 0;rain_draw[38][81] = 0;rain_draw[39][81] = 0;rain_draw[40][81] = 0;rain_draw[41][81] = 0;rain_draw[42][81] = 0;rain_draw[43][81] = 0;rain_draw[44][81] = 0;rain_draw[45][81] = 0;rain_draw[46][81] = 0;rain_draw[47][81] = 0;rain_draw[48][81] = 0;rain_draw[49][81] = 0;rain_draw[50][81] = 0;rain_draw[51][81] = 0;rain_draw[52][81] = 0;rain_draw[53][81] = 0;rain_draw[54][81] = 0;rain_draw[55][81] = 0;rain_draw[56][81] = 0;rain_draw[57][81] = 0;rain_draw[58][81] = 0;rain_draw[59][81] = 0;rain_draw[60][81] = 0;rain_draw[61][81] = 0;rain_draw[62][81] = 1;rain_draw[63][81] = 1;rain_draw[64][81] = 1;rain_draw[65][81] = 0;rain_draw[66][81] = 0;rain_draw[67][81] = 0;rain_draw[68][81] = 0;rain_draw[69][81] = 0;rain_draw[70][81] = 0;rain_draw[71][81] = 0;rain_draw[72][81] = 0;rain_draw[73][81] = 0;rain_draw[74][81] = 0;rain_draw[75][81] = 0;rain_draw[76][81] = 0;rain_draw[77][81] = 0;rain_draw[78][81] = 0;rain_draw[79][81] = 0;rain_draw[80][81] = 0;rain_draw[81][81] = 0;rain_draw[82][81] = 0;rain_draw[83][81] = 0;rain_draw[84][81] = 0;rain_draw[85][81] = 0;rain_draw[86][81] = 0;rain_draw[87][81] = 0;rain_draw[88][81] = 0;rain_draw[89][81] = 0;rain_draw[90][81] = 0;rain_draw[91][81] = 0;rain_draw[92][81] = 0;rain_draw[93][81] = 0;rain_draw[94][81] = 0;rain_draw[95][81] = 0;
        rain_draw[0][82] = 0;rain_draw[1][82] = 0;rain_draw[2][82] = 0;rain_draw[3][82] = 0;rain_draw[4][82] = 0;rain_draw[5][82] = 0;rain_draw[6][82] = 0;rain_draw[7][82] = 0;rain_draw[8][82] = 0;rain_draw[9][82] = 0;rain_draw[10][82] = 0;rain_draw[11][82] = 0;rain_draw[12][82] = 0;rain_draw[13][82] = 0;rain_draw[14][82] = 0;rain_draw[15][82] = 0;rain_draw[16][82] = 0;rain_draw[17][82] = 0;rain_draw[18][82] = 0;rain_draw[19][82] = 0;rain_draw[20][82] = 0;rain_draw[21][82] = 0;rain_draw[22][82] = 0;rain_draw[23][82] = 0;rain_draw[24][82] = 0;rain_draw[25][82] = 0;rain_draw[26][82] = 0;rain_draw[27][82] = 1;rain_draw[28][82] = 1;rain_draw[29][82] = 1;rain_draw[30][82] = 0;rain_draw[31][82] = 0;rain_draw[32][82] = 0;rain_draw[33][82] = 0;rain_draw[34][82] = 0;rain_draw[35][82] = 0;rain_draw[36][82] = 0;rain_draw[37][82] = 0;rain_draw[38][82] = 0;rain_draw[39][82] = 0;rain_draw[40][82] = 0;rain_draw[41][82] = 0;rain_draw[42][82] = 0;rain_draw[43][82] = 0;rain_draw[44][82] = 0;rain_draw[45][82] = 0;rain_draw[46][82] = 0;rain_draw[47][82] = 0;rain_draw[48][82] = 0;rain_draw[49][82] = 0;rain_draw[50][82] = 0;rain_draw[51][82] = 0;rain_draw[52][82] = 0;rain_draw[53][82] = 0;rain_draw[54][82] = 0;rain_draw[55][82] = 0;rain_draw[56][82] = 0;rain_draw[57][82] = 0;rain_draw[58][82] = 0;rain_draw[59][82] = 0;rain_draw[60][82] = 0;rain_draw[61][82] = 0;rain_draw[62][82] = 0;rain_draw[63][82] = 0;rain_draw[64][82] = 0;rain_draw[65][82] = 0;rain_draw[66][82] = 0;rain_draw[67][82] = 0;rain_draw[68][82] = 0;rain_draw[69][82] = 0;rain_draw[70][82] = 0;rain_draw[71][82] = 0;rain_draw[72][82] = 0;rain_draw[73][82] = 0;rain_draw[74][82] = 0;rain_draw[75][82] = 0;rain_draw[76][82] = 0;rain_draw[77][82] = 0;rain_draw[78][82] = 0;rain_draw[79][82] = 0;rain_draw[80][82] = 0;rain_draw[81][82] = 0;rain_draw[82][82] = 0;rain_draw[83][82] = 0;rain_draw[84][82] = 0;rain_draw[85][82] = 0;rain_draw[86][82] = 0;rain_draw[87][82] = 0;rain_draw[88][82] = 0;rain_draw[89][82] = 0;rain_draw[90][82] = 0;rain_draw[91][82] = 0;rain_draw[92][82] = 0;rain_draw[93][82] = 0;rain_draw[94][82] = 0;rain_draw[95][82] = 0;
        rain_draw[0][83] = 0;rain_draw[1][83] = 0;rain_draw[2][83] = 0;rain_draw[3][83] = 0;rain_draw[4][83] = 0;rain_draw[5][83] = 0;rain_draw[6][83] = 0;rain_draw[7][83] = 0;rain_draw[8][83] = 0;rain_draw[9][83] = 0;rain_draw[10][83] = 0;rain_draw[11][83] = 0;rain_draw[12][83] = 0;rain_draw[13][83] = 0;rain_draw[14][83] = 0;rain_draw[15][83] = 0;rain_draw[16][83] = 0;rain_draw[17][83] = 0;rain_draw[18][83] = 0;rain_draw[19][83] = 0;rain_draw[20][83] = 0;rain_draw[21][83] = 0;rain_draw[22][83] = 0;rain_draw[23][83] = 0;rain_draw[24][83] = 0;rain_draw[25][83] = 0;rain_draw[26][83] = 1;rain_draw[27][83] = 1;rain_draw[28][83] = 1;rain_draw[29][83] = 0;rain_draw[30][83] = 0;rain_draw[31][83] = 0;rain_draw[32][83] = 0;rain_draw[33][83] = 0;rain_draw[34][83] = 0;rain_draw[35][83] = 0;rain_draw[36][83] = 0;rain_draw[37][83] = 0;rain_draw[38][83] = 0;rain_draw[39][83] = 0;rain_draw[40][83] = 0;rain_draw[41][83] = 0;rain_draw[42][83] = 0;rain_draw[43][83] = 0;rain_draw[44][83] = 0;rain_draw[45][83] = 0;rain_draw[46][83] = 0;rain_draw[47][83] = 0;rain_draw[48][83] = 0;rain_draw[49][83] = 0;rain_draw[50][83] = 0;rain_draw[51][83] = 0;rain_draw[52][83] = 0;rain_draw[53][83] = 0;rain_draw[54][83] = 0;rain_draw[55][83] = 0;rain_draw[56][83] = 0;rain_draw[57][83] = 0;rain_draw[58][83] = 0;rain_draw[59][83] = 0;rain_draw[60][83] = 0;rain_draw[61][83] = 0;rain_draw[62][83] = 0;rain_draw[63][83] = 0;rain_draw[64][83] = 0;rain_draw[65][83] = 0;rain_draw[66][83] = 0;rain_draw[67][83] = 0;rain_draw[68][83] = 0;rain_draw[69][83] = 0;rain_draw[70][83] = 0;rain_draw[71][83] = 0;rain_draw[72][83] = 0;rain_draw[73][83] = 0;rain_draw[74][83] = 0;rain_draw[75][83] = 0;rain_draw[76][83] = 0;rain_draw[77][83] = 0;rain_draw[78][83] = 0;rain_draw[79][83] = 0;rain_draw[80][83] = 0;rain_draw[81][83] = 0;rain_draw[82][83] = 0;rain_draw[83][83] = 0;rain_draw[84][83] = 0;rain_draw[85][83] = 0;rain_draw[86][83] = 0;rain_draw[87][83] = 0;rain_draw[88][83] = 0;rain_draw[89][83] = 0;rain_draw[90][83] = 0;rain_draw[91][83] = 0;rain_draw[92][83] = 0;rain_draw[93][83] = 0;rain_draw[94][83] = 0;rain_draw[95][83] = 0;
        rain_draw[0][84] = 0;rain_draw[1][84] = 0;rain_draw[2][84] = 0;rain_draw[3][84] = 0;rain_draw[4][84] = 0;rain_draw[5][84] = 0;rain_draw[6][84] = 0;rain_draw[7][84] = 0;rain_draw[8][84] = 0;rain_draw[9][84] = 0;rain_draw[10][84] = 0;rain_draw[11][84] = 0;rain_draw[12][84] = 0;rain_draw[13][84] = 0;rain_draw[14][84] = 0;rain_draw[15][84] = 0;rain_draw[16][84] = 0;rain_draw[17][84] = 0;rain_draw[18][84] = 0;rain_draw[19][84] = 0;rain_draw[20][84] = 0;rain_draw[21][84] = 0;rain_draw[22][84] = 0;rain_draw[23][84] = 0;rain_draw[24][84] = 0;rain_draw[25][84] = 1;rain_draw[26][84] = 1;rain_draw[27][84] = 1;rain_draw[28][84] = 0;rain_draw[29][84] = 0;rain_draw[30][84] = 0;rain_draw[31][84] = 0;rain_draw[32][84] = 0;rain_draw[33][84] = 0;rain_draw[34][84] = 0;rain_draw[35][84] = 0;rain_draw[36][84] = 0;rain_draw[37][84] = 0;rain_draw[38][84] = 0;rain_draw[39][84] = 0;rain_draw[40][84] = 0;rain_draw[41][84] = 0;rain_draw[42][84] = 0;rain_draw[43][84] = 0;rain_draw[44][84] = 0;rain_draw[45][84] = 0;rain_draw[46][84] = 0;rain_draw[47][84] = 0;rain_draw[48][84] = 0;rain_draw[49][84] = 0;rain_draw[50][84] = 0;rain_draw[51][84] = 0;rain_draw[52][84] = 0;rain_draw[53][84] = 0;rain_draw[54][84] = 0;rain_draw[55][84] = 0;rain_draw[56][84] = 0;rain_draw[57][84] = 0;rain_draw[58][84] = 0;rain_draw[59][84] = 0;rain_draw[60][84] = 0;rain_draw[61][84] = 0;rain_draw[62][84] = 0;rain_draw[63][84] = 0;rain_draw[64][84] = 0;rain_draw[65][84] = 0;rain_draw[66][84] = 0;rain_draw[67][84] = 0;rain_draw[68][84] = 0;rain_draw[69][84] = 0;rain_draw[70][84] = 0;rain_draw[71][84] = 0;rain_draw[72][84] = 0;rain_draw[73][84] = 0;rain_draw[74][84] = 0;rain_draw[75][84] = 0;rain_draw[76][84] = 0;rain_draw[77][84] = 0;rain_draw[78][84] = 0;rain_draw[79][84] = 0;rain_draw[80][84] = 0;rain_draw[81][84] = 0;rain_draw[82][84] = 0;rain_draw[83][84] = 0;rain_draw[84][84] = 0;rain_draw[85][84] = 1;rain_draw[86][84] = 1;rain_draw[87][84] = 1;rain_draw[88][84] = 0;rain_draw[89][84] = 0;rain_draw[90][84] = 0;rain_draw[91][84] = 0;rain_draw[92][84] = 0;rain_draw[93][84] = 0;rain_draw[94][84] = 0;rain_draw[95][84] = 0;
        rain_draw[0][85] = 0;rain_draw[1][85] = 0;rain_draw[2][85] = 0;rain_draw[3][85] = 0;rain_draw[4][85] = 0;rain_draw[5][85] = 0;rain_draw[6][85] = 0;rain_draw[7][85] = 0;rain_draw[8][85] = 0;rain_draw[9][85] = 0;rain_draw[10][85] = 0;rain_draw[11][85] = 0;rain_draw[12][85] = 0;rain_draw[13][85] = 0;rain_draw[14][85] = 0;rain_draw[15][85] = 0;rain_draw[16][85] = 0;rain_draw[17][85] = 0;rain_draw[18][85] = 0;rain_draw[19][85] = 0;rain_draw[20][85] = 0;rain_draw[21][85] = 0;rain_draw[22][85] = 0;rain_draw[23][85] = 0;rain_draw[24][85] = 1;rain_draw[25][85] = 1;rain_draw[26][85] = 1;rain_draw[27][85] = 0;rain_draw[28][85] = 0;rain_draw[29][85] = 0;rain_draw[30][85] = 0;rain_draw[31][85] = 0;rain_draw[32][85] = 0;rain_draw[33][85] = 0;rain_draw[34][85] = 0;rain_draw[35][85] = 0;rain_draw[36][85] = 0;rain_draw[37][85] = 0;rain_draw[38][85] = 0;rain_draw[39][85] = 0;rain_draw[40][85] = 0;rain_draw[41][85] = 0;rain_draw[42][85] = 0;rain_draw[43][85] = 0;rain_draw[44][85] = 0;rain_draw[45][85] = 0;rain_draw[46][85] = 0;rain_draw[47][85] = 0;rain_draw[48][85] = 0;rain_draw[49][85] = 0;rain_draw[50][85] = 0;rain_draw[51][85] = 0;rain_draw[52][85] = 0;rain_draw[53][85] = 0;rain_draw[54][85] = 0;rain_draw[55][85] = 0;rain_draw[56][85] = 0;rain_draw[57][85] = 0;rain_draw[58][85] = 0;rain_draw[59][85] = 0;rain_draw[60][85] = 0;rain_draw[61][85] = 0;rain_draw[62][85] = 0;rain_draw[63][85] = 0;rain_draw[64][85] = 0;rain_draw[65][85] = 0;rain_draw[66][85] = 0;rain_draw[67][85] = 0;rain_draw[68][85] = 0;rain_draw[69][85] = 0;rain_draw[70][85] = 0;rain_draw[71][85] = 0;rain_draw[72][85] = 0;rain_draw[73][85] = 0;rain_draw[74][85] = 0;rain_draw[75][85] = 0;rain_draw[76][85] = 0;rain_draw[77][85] = 0;rain_draw[78][85] = 0;rain_draw[79][85] = 0;rain_draw[80][85] = 0;rain_draw[81][85] = 0;rain_draw[82][85] = 0;rain_draw[83][85] = 0;rain_draw[84][85] = 1;rain_draw[85][85] = 1;rain_draw[86][85] = 1;rain_draw[87][85] = 0;rain_draw[88][85] = 0;rain_draw[89][85] = 0;rain_draw[90][85] = 0;rain_draw[91][85] = 0;rain_draw[92][85] = 0;rain_draw[93][85] = 0;rain_draw[94][85] = 0;rain_draw[95][85] = 0;
        rain_draw[0][86] = 0;rain_draw[1][86] = 0;rain_draw[2][86] = 0;rain_draw[3][86] = 0;rain_draw[4][86] = 0;rain_draw[5][86] = 0;rain_draw[6][86] = 0;rain_draw[7][86] = 0;rain_draw[8][86] = 0;rain_draw[9][86] = 0;rain_draw[10][86] = 0;rain_draw[11][86] = 0;rain_draw[12][86] = 0;rain_draw[13][86] = 0;rain_draw[14][86] = 0;rain_draw[15][86] = 0;rain_draw[16][86] = 0;rain_draw[17][86] = 0;rain_draw[18][86] = 0;rain_draw[19][86] = 0;rain_draw[20][86] = 0;rain_draw[21][86] = 0;rain_draw[22][86] = 0;rain_draw[23][86] = 1;rain_draw[24][86] = 1;rain_draw[25][86] = 1;rain_draw[26][86] = 0;rain_draw[27][86] = 0;rain_draw[28][86] = 0;rain_draw[29][86] = 0;rain_draw[30][86] = 0;rain_draw[31][86] = 0;rain_draw[32][86] = 0;rain_draw[33][86] = 0;rain_draw[34][86] = 0;rain_draw[35][86] = 0;rain_draw[36][86] = 0;rain_draw[37][86] = 0;rain_draw[38][86] = 0;rain_draw[39][86] = 0;rain_draw[40][86] = 0;rain_draw[41][86] = 0;rain_draw[42][86] = 0;rain_draw[43][86] = 0;rain_draw[44][86] = 0;rain_draw[45][86] = 0;rain_draw[46][86] = 0;rain_draw[47][86] = 0;rain_draw[48][86] = 0;rain_draw[49][86] = 0;rain_draw[50][86] = 0;rain_draw[51][86] = 0;rain_draw[52][86] = 0;rain_draw[53][86] = 0;rain_draw[54][86] = 0;rain_draw[55][86] = 0;rain_draw[56][86] = 0;rain_draw[57][86] = 0;rain_draw[58][86] = 0;rain_draw[59][86] = 0;rain_draw[60][86] = 0;rain_draw[61][86] = 0;rain_draw[62][86] = 0;rain_draw[63][86] = 0;rain_draw[64][86] = 0;rain_draw[65][86] = 0;rain_draw[66][86] = 0;rain_draw[67][86] = 0;rain_draw[68][86] = 0;rain_draw[69][86] = 0;rain_draw[70][86] = 0;rain_draw[71][86] = 0;rain_draw[72][86] = 0;rain_draw[73][86] = 0;rain_draw[74][86] = 0;rain_draw[75][86] = 0;rain_draw[76][86] = 0;rain_draw[77][86] = 0;rain_draw[78][86] = 0;rain_draw[79][86] = 0;rain_draw[80][86] = 0;rain_draw[81][86] = 0;rain_draw[82][86] = 0;rain_draw[83][86] = 1;rain_draw[84][86] = 1;rain_draw[85][86] = 1;rain_draw[86][86] = 0;rain_draw[87][86] = 0;rain_draw[88][86] = 0;rain_draw[89][86] = 0;rain_draw[90][86] = 0;rain_draw[91][86] = 0;rain_draw[92][86] = 0;rain_draw[93][86] = 0;rain_draw[94][86] = 0;rain_draw[95][86] = 0;
        rain_draw[0][87] = 0;rain_draw[1][87] = 0;rain_draw[2][87] = 0;rain_draw[3][87] = 0;rain_draw[4][87] = 0;rain_draw[5][87] = 0;rain_draw[6][87] = 0;rain_draw[7][87] = 0;rain_draw[8][87] = 0;rain_draw[9][87] = 0;rain_draw[10][87] = 0;rain_draw[11][87] = 0;rain_draw[12][87] = 0;rain_draw[13][87] = 0;rain_draw[14][87] = 0;rain_draw[15][87] = 0;rain_draw[16][87] = 0;rain_draw[17][87] = 0;rain_draw[18][87] = 0;rain_draw[19][87] = 0;rain_draw[20][87] = 0;rain_draw[21][87] = 0;rain_draw[22][87] = 0;rain_draw[23][87] = 0;rain_draw[24][87] = 0;rain_draw[25][87] = 0;rain_draw[26][87] = 0;rain_draw[27][87] = 0;rain_draw[28][87] = 0;rain_draw[29][87] = 0;rain_draw[30][87] = 0;rain_draw[31][87] = 0;rain_draw[32][87] = 0;rain_draw[33][87] = 0;rain_draw[34][87] = 0;rain_draw[35][87] = 0;rain_draw[36][87] = 0;rain_draw[37][87] = 0;rain_draw[38][87] = 0;rain_draw[39][87] = 0;rain_draw[40][87] = 0;rain_draw[41][87] = 0;rain_draw[42][87] = 0;rain_draw[43][87] = 0;rain_draw[44][87] = 0;rain_draw[45][87] = 0;rain_draw[46][87] = 0;rain_draw[47][87] = 0;rain_draw[48][87] = 0;rain_draw[49][87] = 0;rain_draw[50][87] = 0;rain_draw[51][87] = 0;rain_draw[52][87] = 0;rain_draw[53][87] = 0;rain_draw[54][87] = 0;rain_draw[55][87] = 0;rain_draw[56][87] = 0;rain_draw[57][87] = 0;rain_draw[58][87] = 0;rain_draw[59][87] = 0;rain_draw[60][87] = 0;rain_draw[61][87] = 0;rain_draw[62][87] = 0;rain_draw[63][87] = 0;rain_draw[64][87] = 0;rain_draw[65][87] = 0;rain_draw[66][87] = 0;rain_draw[67][87] = 0;rain_draw[68][87] = 0;rain_draw[69][87] = 0;rain_draw[70][87] = 0;rain_draw[71][87] = 0;rain_draw[72][87] = 0;rain_draw[73][87] = 0;rain_draw[74][87] = 0;rain_draw[75][87] = 0;rain_draw[76][87] = 0;rain_draw[77][87] = 0;rain_draw[78][87] = 0;rain_draw[79][87] = 0;rain_draw[80][87] = 0;rain_draw[81][87] = 0;rain_draw[82][87] = 1;rain_draw[83][87] = 1;rain_draw[84][87] = 1;rain_draw[85][87] = 0;rain_draw[86][87] = 0;rain_draw[87][87] = 0;rain_draw[88][87] = 0;rain_draw[89][87] = 0;rain_draw[90][87] = 0;rain_draw[91][87] = 0;rain_draw[92][87] = 0;rain_draw[93][87] = 0;rain_draw[94][87] = 0;rain_draw[95][87] = 0;
        rain_draw[0][88] = 0;rain_draw[1][88] = 0;rain_draw[2][88] = 0;rain_draw[3][88] = 0;rain_draw[4][88] = 0;rain_draw[5][88] = 0;rain_draw[6][88] = 0;rain_draw[7][88] = 0;rain_draw[8][88] = 0;rain_draw[9][88] = 0;rain_draw[10][88] = 0;rain_draw[11][88] = 0;rain_draw[12][88] = 0;rain_draw[13][88] = 0;rain_draw[14][88] = 0;rain_draw[15][88] = 0;rain_draw[16][88] = 0;rain_draw[17][88] = 0;rain_draw[18][88] = 0;rain_draw[19][88] = 0;rain_draw[20][88] = 0;rain_draw[21][88] = 0;rain_draw[22][88] = 0;rain_draw[23][88] = 0;rain_draw[24][88] = 0;rain_draw[25][88] = 0;rain_draw[26][88] = 0;rain_draw[27][88] = 0;rain_draw[28][88] = 0;rain_draw[29][88] = 0;rain_draw[30][88] = 0;rain_draw[31][88] = 0;rain_draw[32][88] = 0;rain_draw[33][88] = 0;rain_draw[34][88] = 0;rain_draw[35][88] = 0;rain_draw[36][88] = 0;rain_draw[37][88] = 0;rain_draw[38][88] = 0;rain_draw[39][88] = 0;rain_draw[40][88] = 0;rain_draw[41][88] = 0;rain_draw[42][88] = 0;rain_draw[43][88] = 0;rain_draw[44][88] = 0;rain_draw[45][88] = 0;rain_draw[46][88] = 0;rain_draw[47][88] = 0;rain_draw[48][88] = 0;rain_draw[49][88] = 0;rain_draw[50][88] = 0;rain_draw[51][88] = 0;rain_draw[52][88] = 0;rain_draw[53][88] = 0;rain_draw[54][88] = 0;rain_draw[55][88] = 0;rain_draw[56][88] = 0;rain_draw[57][88] = 0;rain_draw[58][88] = 0;rain_draw[59][88] = 0;rain_draw[60][88] = 0;rain_draw[61][88] = 0;rain_draw[62][88] = 0;rain_draw[63][88] = 0;rain_draw[64][88] = 0;rain_draw[65][88] = 0;rain_draw[66][88] = 0;rain_draw[67][88] = 0;rain_draw[68][88] = 0;rain_draw[69][88] = 0;rain_draw[70][88] = 0;rain_draw[71][88] = 0;rain_draw[72][88] = 0;rain_draw[73][88] = 0;rain_draw[74][88] = 0;rain_draw[75][88] = 0;rain_draw[76][88] = 0;rain_draw[77][88] = 0;rain_draw[78][88] = 0;rain_draw[79][88] = 0;rain_draw[80][88] = 0;rain_draw[81][88] = 1;rain_draw[82][88] = 1;rain_draw[83][88] = 1;rain_draw[84][88] = 0;rain_draw[85][88] = 0;rain_draw[86][88] = 0;rain_draw[87][88] = 0;rain_draw[88][88] = 0;rain_draw[89][88] = 0;rain_draw[90][88] = 0;rain_draw[91][88] = 0;rain_draw[92][88] = 0;rain_draw[93][88] = 0;rain_draw[94][88] = 0;rain_draw[95][88] = 0;
        rain_draw[0][89] = 0;rain_draw[1][89] = 0;rain_draw[2][89] = 0;rain_draw[3][89] = 0;rain_draw[4][89] = 0;rain_draw[5][89] = 0;rain_draw[6][89] = 0;rain_draw[7][89] = 0;rain_draw[8][89] = 0;rain_draw[9][89] = 0;rain_draw[10][89] = 0;rain_draw[11][89] = 0;rain_draw[12][89] = 0;rain_draw[13][89] = 0;rain_draw[14][89] = 0;rain_draw[15][89] = 0;rain_draw[16][89] = 0;rain_draw[17][89] = 0;rain_draw[18][89] = 0;rain_draw[19][89] = 0;rain_draw[20][89] = 0;rain_draw[21][89] = 0;rain_draw[22][89] = 0;rain_draw[23][89] = 0;rain_draw[24][89] = 0;rain_draw[25][89] = 0;rain_draw[26][89] = 0;rain_draw[27][89] = 0;rain_draw[28][89] = 0;rain_draw[29][89] = 0;rain_draw[30][89] = 0;rain_draw[31][89] = 0;rain_draw[32][89] = 0;rain_draw[33][89] = 0;rain_draw[34][89] = 0;rain_draw[35][89] = 0;rain_draw[36][89] = 0;rain_draw[37][89] = 0;rain_draw[38][89] = 0;rain_draw[39][89] = 0;rain_draw[40][89] = 0;rain_draw[41][89] = 0;rain_draw[42][89] = 0;rain_draw[43][89] = 0;rain_draw[44][89] = 0;rain_draw[45][89] = 0;rain_draw[46][89] = 0;rain_draw[47][89] = 0;rain_draw[48][89] = 0;rain_draw[49][89] = 0;rain_draw[50][89] = 0;rain_draw[51][89] = 0;rain_draw[52][89] = 1;rain_draw[53][89] = 1;rain_draw[54][89] = 1;rain_draw[55][89] = 0;rain_draw[56][89] = 0;rain_draw[57][89] = 0;rain_draw[58][89] = 0;rain_draw[59][89] = 0;rain_draw[60][89] = 0;rain_draw[61][89] = 0;rain_draw[62][89] = 0;rain_draw[63][89] = 0;rain_draw[64][89] = 0;rain_draw[65][89] = 0;rain_draw[66][89] = 0;rain_draw[67][89] = 0;rain_draw[68][89] = 0;rain_draw[69][89] = 0;rain_draw[70][89] = 0;rain_draw[71][89] = 0;rain_draw[72][89] = 0;rain_draw[73][89] = 0;rain_draw[74][89] = 0;rain_draw[75][89] = 0;rain_draw[76][89] = 0;rain_draw[77][89] = 0;rain_draw[78][89] = 0;rain_draw[79][89] = 0;rain_draw[80][89] = 1;rain_draw[81][89] = 1;rain_draw[82][89] = 1;rain_draw[83][89] = 0;rain_draw[84][89] = 0;rain_draw[85][89] = 0;rain_draw[86][89] = 0;rain_draw[87][89] = 0;rain_draw[88][89] = 0;rain_draw[89][89] = 0;rain_draw[90][89] = 0;rain_draw[91][89] = 0;rain_draw[92][89] = 0;rain_draw[93][89] = 0;rain_draw[94][89] = 0;rain_draw[95][89] = 0;
        rain_draw[0][90] = 0;rain_draw[1][90] = 0;rain_draw[2][90] = 0;rain_draw[3][90] = 0;rain_draw[4][90] = 0;rain_draw[5][90] = 0;rain_draw[6][90] = 0;rain_draw[7][90] = 0;rain_draw[8][90] = 0;rain_draw[9][90] = 0;rain_draw[10][90] = 0;rain_draw[11][90] = 0;rain_draw[12][90] = 0;rain_draw[13][90] = 0;rain_draw[14][90] = 0;rain_draw[15][90] = 0;rain_draw[16][90] = 0;rain_draw[17][90] = 0;rain_draw[18][90] = 0;rain_draw[19][90] = 0;rain_draw[20][90] = 0;rain_draw[21][90] = 0;rain_draw[22][90] = 0;rain_draw[23][90] = 0;rain_draw[24][90] = 0;rain_draw[25][90] = 0;rain_draw[26][90] = 0;rain_draw[27][90] = 0;rain_draw[28][90] = 0;rain_draw[29][90] = 0;rain_draw[30][90] = 0;rain_draw[31][90] = 0;rain_draw[32][90] = 0;rain_draw[33][90] = 0;rain_draw[34][90] = 0;rain_draw[35][90] = 0;rain_draw[36][90] = 0;rain_draw[37][90] = 0;rain_draw[38][90] = 0;rain_draw[39][90] = 0;rain_draw[40][90] = 0;rain_draw[41][90] = 0;rain_draw[42][90] = 0;rain_draw[43][90] = 0;rain_draw[44][90] = 0;rain_draw[45][90] = 0;rain_draw[46][90] = 0;rain_draw[47][90] = 0;rain_draw[48][90] = 0;rain_draw[49][90] = 0;rain_draw[50][90] = 0;rain_draw[51][90] = 1;rain_draw[52][90] = 1;rain_draw[53][90] = 1;rain_draw[54][90] = 0;rain_draw[55][90] = 0;rain_draw[56][90] = 0;rain_draw[57][90] = 0;rain_draw[58][90] = 0;rain_draw[59][90] = 0;rain_draw[60][90] = 0;rain_draw[61][90] = 0;rain_draw[62][90] = 0;rain_draw[63][90] = 0;rain_draw[64][90] = 0;rain_draw[65][90] = 0;rain_draw[66][90] = 0;rain_draw[67][90] = 0;rain_draw[68][90] = 0;rain_draw[69][90] = 0;rain_draw[70][90] = 0;rain_draw[71][90] = 0;rain_draw[72][90] = 0;rain_draw[73][90] = 0;rain_draw[74][90] = 0;rain_draw[75][90] = 0;rain_draw[76][90] = 0;rain_draw[77][90] = 0;rain_draw[78][90] = 0;rain_draw[79][90] = 1;rain_draw[80][90] = 1;rain_draw[81][90] = 1;rain_draw[82][90] = 0;rain_draw[83][90] = 0;rain_draw[84][90] = 0;rain_draw[85][90] = 0;rain_draw[86][90] = 0;rain_draw[87][90] = 0;rain_draw[88][90] = 0;rain_draw[89][90] = 0;rain_draw[90][90] = 0;rain_draw[91][90] = 0;rain_draw[92][90] = 0;rain_draw[93][90] = 0;rain_draw[94][90] = 0;rain_draw[95][90] = 0;
        rain_draw[0][91] = 0;rain_draw[1][91] = 0;rain_draw[2][91] = 0;rain_draw[3][91] = 0;rain_draw[4][91] = 0;rain_draw[5][91] = 0;rain_draw[6][91] = 0;rain_draw[7][91] = 0;rain_draw[8][91] = 0;rain_draw[9][91] = 0;rain_draw[10][91] = 0;rain_draw[11][91] = 0;rain_draw[12][91] = 0;rain_draw[13][91] = 0;rain_draw[14][91] = 0;rain_draw[15][91] = 0;rain_draw[16][91] = 0;rain_draw[17][91] = 0;rain_draw[18][91] = 0;rain_draw[19][91] = 0;rain_draw[20][91] = 0;rain_draw[21][91] = 0;rain_draw[22][91] = 0;rain_draw[23][91] = 0;rain_draw[24][91] = 0;rain_draw[25][91] = 0;rain_draw[26][91] = 0;rain_draw[27][91] = 0;rain_draw[28][91] = 0;rain_draw[29][91] = 0;rain_draw[30][91] = 0;rain_draw[31][91] = 0;rain_draw[32][91] = 0;rain_draw[33][91] = 0;rain_draw[34][91] = 0;rain_draw[35][91] = 0;rain_draw[36][91] = 0;rain_draw[37][91] = 0;rain_draw[38][91] = 0;rain_draw[39][91] = 0;rain_draw[40][91] = 0;rain_draw[41][91] = 0;rain_draw[42][91] = 0;rain_draw[43][91] = 0;rain_draw[44][91] = 0;rain_draw[45][91] = 0;rain_draw[46][91] = 0;rain_draw[47][91] = 0;rain_draw[48][91] = 0;rain_draw[49][91] = 0;rain_draw[50][91] = 1;rain_draw[51][91] = 1;rain_draw[52][91] = 1;rain_draw[53][91] = 0;rain_draw[54][91] = 0;rain_draw[55][91] = 0;rain_draw[56][91] = 0;rain_draw[57][91] = 0;rain_draw[58][91] = 0;rain_draw[59][91] = 0;rain_draw[60][91] = 0;rain_draw[61][91] = 0;rain_draw[62][91] = 0;rain_draw[63][91] = 0;rain_draw[64][91] = 0;rain_draw[65][91] = 0;rain_draw[66][91] = 0;rain_draw[67][91] = 0;rain_draw[68][91] = 0;rain_draw[69][91] = 0;rain_draw[70][91] = 0;rain_draw[71][91] = 0;rain_draw[72][91] = 0;rain_draw[73][91] = 0;rain_draw[74][91] = 0;rain_draw[75][91] = 0;rain_draw[76][91] = 0;rain_draw[77][91] = 0;rain_draw[78][91] = 0;rain_draw[79][91] = 0;rain_draw[80][91] = 0;rain_draw[81][91] = 0;rain_draw[82][91] = 0;rain_draw[83][91] = 0;rain_draw[84][91] = 0;rain_draw[85][91] = 0;rain_draw[86][91] = 0;rain_draw[87][91] = 0;rain_draw[88][91] = 0;rain_draw[89][91] = 0;rain_draw[90][91] = 0;rain_draw[91][91] = 0;rain_draw[92][91] = 0;rain_draw[93][91] = 0;rain_draw[94][91] = 0;rain_draw[95][91] = 0;
        rain_draw[0][92] = 0;rain_draw[1][92] = 0;rain_draw[2][92] = 0;rain_draw[3][92] = 0;rain_draw[4][92] = 0;rain_draw[5][92] = 0;rain_draw[6][92] = 0;rain_draw[7][92] = 0;rain_draw[8][92] = 0;rain_draw[9][92] = 0;rain_draw[10][92] = 0;rain_draw[11][92] = 0;rain_draw[12][92] = 0;rain_draw[13][92] = 0;rain_draw[14][92] = 0;rain_draw[15][92] = 0;rain_draw[16][92] = 0;rain_draw[17][92] = 0;rain_draw[18][92] = 0;rain_draw[19][92] = 0;rain_draw[20][92] = 0;rain_draw[21][92] = 0;rain_draw[22][92] = 0;rain_draw[23][92] = 0;rain_draw[24][92] = 0;rain_draw[25][92] = 0;rain_draw[26][92] = 0;rain_draw[27][92] = 0;rain_draw[28][92] = 0;rain_draw[29][92] = 0;rain_draw[30][92] = 0;rain_draw[31][92] = 0;rain_draw[32][92] = 0;rain_draw[33][92] = 0;rain_draw[34][92] = 0;rain_draw[35][92] = 0;rain_draw[36][92] = 0;rain_draw[37][92] = 0;rain_draw[38][92] = 0;rain_draw[39][92] = 0;rain_draw[40][92] = 0;rain_draw[41][92] = 0;rain_draw[42][92] = 0;rain_draw[43][92] = 0;rain_draw[44][92] = 0;rain_draw[45][92] = 0;rain_draw[46][92] = 0;rain_draw[47][92] = 0;rain_draw[48][92] = 0;rain_draw[49][92] = 1;rain_draw[50][92] = 1;rain_draw[51][92] = 1;rain_draw[52][92] = 0;rain_draw[53][92] = 0;rain_draw[54][92] = 0;rain_draw[55][92] = 0;rain_draw[56][92] = 0;rain_draw[57][92] = 0;rain_draw[58][92] = 0;rain_draw[59][92] = 0;rain_draw[60][92] = 0;rain_draw[61][92] = 0;rain_draw[62][92] = 0;rain_draw[63][92] = 0;rain_draw[64][92] = 0;rain_draw[65][92] = 0;rain_draw[66][92] = 0;rain_draw[67][92] = 0;rain_draw[68][92] = 0;rain_draw[69][92] = 0;rain_draw[70][92] = 0;rain_draw[71][92] = 0;rain_draw[72][92] = 0;rain_draw[73][92] = 0;rain_draw[74][92] = 0;rain_draw[75][92] = 0;rain_draw[76][92] = 0;rain_draw[77][92] = 0;rain_draw[78][92] = 0;rain_draw[79][92] = 0;rain_draw[80][92] = 0;rain_draw[81][92] = 0;rain_draw[82][92] = 0;rain_draw[83][92] = 0;rain_draw[84][92] = 0;rain_draw[85][92] = 0;rain_draw[86][92] = 0;rain_draw[87][92] = 0;rain_draw[88][92] = 0;rain_draw[89][92] = 0;rain_draw[90][92] = 0;rain_draw[91][92] = 0;rain_draw[92][92] = 0;rain_draw[93][92] = 0;rain_draw[94][92] = 0;rain_draw[95][92] = 0;
        rain_draw[0][93] = 0;rain_draw[1][93] = 0;rain_draw[2][93] = 0;rain_draw[3][93] = 0;rain_draw[4][93] = 0;rain_draw[5][93] = 0;rain_draw[6][93] = 0;rain_draw[7][93] = 0;rain_draw[8][93] = 0;rain_draw[9][93] = 0;rain_draw[10][93] = 0;rain_draw[11][93] = 0;rain_draw[12][93] = 0;rain_draw[13][93] = 0;rain_draw[14][93] = 0;rain_draw[15][93] = 0;rain_draw[16][93] = 0;rain_draw[17][93] = 0;rain_draw[18][93] = 0;rain_draw[19][93] = 0;rain_draw[20][93] = 0;rain_draw[21][93] = 0;rain_draw[22][93] = 0;rain_draw[23][93] = 0;rain_draw[24][93] = 0;rain_draw[25][93] = 0;rain_draw[26][93] = 0;rain_draw[27][93] = 0;rain_draw[28][93] = 0;rain_draw[29][93] = 0;rain_draw[30][93] = 0;rain_draw[31][93] = 0;rain_draw[32][93] = 0;rain_draw[33][93] = 0;rain_draw[34][93] = 0;rain_draw[35][93] = 0;rain_draw[36][93] = 0;rain_draw[37][93] = 0;rain_draw[38][93] = 0;rain_draw[39][93] = 0;rain_draw[40][93] = 0;rain_draw[41][93] = 0;rain_draw[42][93] = 0;rain_draw[43][93] = 0;rain_draw[44][93] = 0;rain_draw[45][93] = 0;rain_draw[46][93] = 0;rain_draw[47][93] = 0;rain_draw[48][93] = 1;rain_draw[49][93] = 1;rain_draw[50][93] = 1;rain_draw[51][93] = 0;rain_draw[52][93] = 0;rain_draw[53][93] = 0;rain_draw[54][93] = 0;rain_draw[55][93] = 0;rain_draw[56][93] = 0;rain_draw[57][93] = 0;rain_draw[58][93] = 0;rain_draw[59][93] = 0;rain_draw[60][93] = 0;rain_draw[61][93] = 0;rain_draw[62][93] = 0;rain_draw[63][93] = 0;rain_draw[64][93] = 0;rain_draw[65][93] = 0;rain_draw[66][93] = 0;rain_draw[67][93] = 0;rain_draw[68][93] = 0;rain_draw[69][93] = 0;rain_draw[70][93] = 0;rain_draw[71][93] = 0;rain_draw[72][93] = 0;rain_draw[73][93] = 0;rain_draw[74][93] = 0;rain_draw[75][93] = 0;rain_draw[76][93] = 0;rain_draw[77][93] = 0;rain_draw[78][93] = 0;rain_draw[79][93] = 0;rain_draw[80][93] = 0;rain_draw[81][93] = 0;rain_draw[82][93] = 0;rain_draw[83][93] = 0;rain_draw[84][93] = 0;rain_draw[85][93] = 0;rain_draw[86][93] = 0;rain_draw[87][93] = 0;rain_draw[88][93] = 0;rain_draw[89][93] = 0;rain_draw[90][93] = 0;rain_draw[91][93] = 0;rain_draw[92][93] = 0;rain_draw[93][93] = 0;rain_draw[94][93] = 0;rain_draw[95][93] = 0;
        rain_draw[0][94] = 0;rain_draw[1][94] = 0;rain_draw[2][94] = 0;rain_draw[3][94] = 0;rain_draw[4][94] = 0;rain_draw[5][94] = 0;rain_draw[6][94] = 0;rain_draw[7][94] = 0;rain_draw[8][94] = 0;rain_draw[9][94] = 1;rain_draw[10][94] = 1;rain_draw[11][94] = 1;rain_draw[12][94] = 0;rain_draw[13][94] = 0;rain_draw[14][94] = 0;rain_draw[15][94] = 0;rain_draw[16][94] = 0;rain_draw[17][94] = 0;rain_draw[18][94] = 0;rain_draw[19][94] = 0;rain_draw[20][94] = 0;rain_draw[21][94] = 0;rain_draw[22][94] = 0;rain_draw[23][94] = 0;rain_draw[24][94] = 0;rain_draw[25][94] = 0;rain_draw[26][94] = 0;rain_draw[27][94] = 0;rain_draw[28][94] = 0;rain_draw[29][94] = 0;rain_draw[30][94] = 0;rain_draw[31][94] = 0;rain_draw[32][94] = 0;rain_draw[33][94] = 0;rain_draw[34][94] = 0;rain_draw[35][94] = 0;rain_draw[36][94] = 0;rain_draw[37][94] = 0;rain_draw[38][94] = 0;rain_draw[39][94] = 0;rain_draw[40][94] = 0;rain_draw[41][94] = 0;rain_draw[42][94] = 0;rain_draw[43][94] = 0;rain_draw[44][94] = 0;rain_draw[45][94] = 0;rain_draw[46][94] = 0;rain_draw[47][94] = 1;rain_draw[48][94] = 1;rain_draw[49][94] = 1;rain_draw[50][94] = 0;rain_draw[51][94] = 0;rain_draw[52][94] = 0;rain_draw[53][94] = 0;rain_draw[54][94] = 0;rain_draw[55][94] = 0;rain_draw[56][94] = 0;rain_draw[57][94] = 0;rain_draw[58][94] = 0;rain_draw[59][94] = 0;rain_draw[60][94] = 0;rain_draw[61][94] = 0;rain_draw[62][94] = 0;rain_draw[63][94] = 0;rain_draw[64][94] = 0;rain_draw[65][94] = 0;rain_draw[66][94] = 0;rain_draw[67][94] = 0;rain_draw[68][94] = 0;rain_draw[69][94] = 0;rain_draw[70][94] = 0;rain_draw[71][94] = 0;rain_draw[72][94] = 0;rain_draw[73][94] = 0;rain_draw[74][94] = 0;rain_draw[75][94] = 0;rain_draw[76][94] = 0;rain_draw[77][94] = 0;rain_draw[78][94] = 0;rain_draw[79][94] = 0;rain_draw[80][94] = 0;rain_draw[81][94] = 0;rain_draw[82][94] = 0;rain_draw[83][94] = 0;rain_draw[84][94] = 0;rain_draw[85][94] = 0;rain_draw[86][94] = 0;rain_draw[87][94] = 0;rain_draw[88][94] = 0;rain_draw[89][94] = 0;rain_draw[90][94] = 0;rain_draw[91][94] = 0;rain_draw[92][94] = 0;rain_draw[93][94] = 0;rain_draw[94][94] = 0;rain_draw[95][94] = 0;
        rain_draw[0][95] = 0;rain_draw[1][95] = 0;rain_draw[2][95] = 0;rain_draw[3][95] = 0;rain_draw[4][95] = 0;rain_draw[5][95] = 0;rain_draw[6][95] = 0;rain_draw[7][95] = 0;rain_draw[8][95] = 1;rain_draw[9][95] = 1;rain_draw[10][95] = 1;rain_draw[11][95] = 0;rain_draw[12][95] = 0;rain_draw[13][95] = 0;rain_draw[14][95] = 0;rain_draw[15][95] = 0;rain_draw[16][95] = 0;rain_draw[17][95] = 0;rain_draw[18][95] = 0;rain_draw[19][95] = 0;rain_draw[20][95] = 0;rain_draw[21][95] = 0;rain_draw[22][95] = 0;rain_draw[23][95] = 0;rain_draw[24][95] = 0;rain_draw[25][95] = 0;rain_draw[26][95] = 0;rain_draw[27][95] = 0;rain_draw[28][95] = 0;rain_draw[29][95] = 0;rain_draw[30][95] = 0;rain_draw[31][95] = 0;rain_draw[32][95] = 0;rain_draw[33][95] = 0;rain_draw[34][95] = 0;rain_draw[35][95] = 0;rain_draw[36][95] = 0;rain_draw[37][95] = 0;rain_draw[38][95] = 0;rain_draw[39][95] = 0;rain_draw[40][95] = 0;rain_draw[41][95] = 0;rain_draw[42][95] = 0;rain_draw[43][95] = 0;rain_draw[44][95] = 0;rain_draw[45][95] = 0;rain_draw[46][95] = 1;rain_draw[47][95] = 1;rain_draw[48][95] = 1;rain_draw[49][95] = 0;rain_draw[50][95] = 0;rain_draw[51][95] = 0;rain_draw[52][95] = 0;rain_draw[53][95] = 0;rain_draw[54][95] = 0;rain_draw[55][95] = 0;rain_draw[56][95] = 0;rain_draw[57][95] = 0;rain_draw[58][95] = 0;rain_draw[59][95] = 0;rain_draw[60][95] = 0;rain_draw[61][95] = 0;rain_draw[62][95] = 0;rain_draw[63][95] = 0;rain_draw[64][95] = 0;rain_draw[65][95] = 0;rain_draw[66][95] = 0;rain_draw[67][95] = 0;rain_draw[68][95] = 0;rain_draw[69][95] = 0;rain_draw[70][95] = 0;rain_draw[71][95] = 0;rain_draw[72][95] = 0;rain_draw[73][95] = 0;rain_draw[74][95] = 0;rain_draw[75][95] = 0;rain_draw[76][95] = 0;rain_draw[77][95] = 0;rain_draw[78][95] = 0;rain_draw[79][95] = 0;rain_draw[80][95] = 0;rain_draw[81][95] = 0;rain_draw[82][95] = 0;rain_draw[83][95] = 0;rain_draw[84][95] = 0;rain_draw[85][95] = 0;rain_draw[86][95] = 0;rain_draw[87][95] = 0;rain_draw[88][95] = 0;rain_draw[89][95] = 0;rain_draw[90][95] = 0;rain_draw[91][95] = 0;rain_draw[92][95] = 0;rain_draw[93][95] = 0;rain_draw[94][95] = 0;rain_draw[95][95] = 0;
        rain_draw[0][96] = 0;rain_draw[1][96] = 0;rain_draw[2][96] = 0;rain_draw[3][96] = 0;rain_draw[4][96] = 0;rain_draw[5][96] = 0;rain_draw[6][96] = 0;rain_draw[7][96] = 1;rain_draw[8][96] = 1;rain_draw[9][96] = 1;rain_draw[10][96] = 0;rain_draw[11][96] = 0;rain_draw[12][96] = 0;rain_draw[13][96] = 0;rain_draw[14][96] = 0;rain_draw[15][96] = 0;rain_draw[16][96] = 0;rain_draw[17][96] = 0;rain_draw[18][96] = 0;rain_draw[19][96] = 0;rain_draw[20][96] = 0;rain_draw[21][96] = 0;rain_draw[22][96] = 0;rain_draw[23][96] = 0;rain_draw[24][96] = 0;rain_draw[25][96] = 0;rain_draw[26][96] = 0;rain_draw[27][96] = 0;rain_draw[28][96] = 0;rain_draw[29][96] = 0;rain_draw[30][96] = 0;rain_draw[31][96] = 0;rain_draw[32][96] = 0;rain_draw[33][96] = 0;rain_draw[34][96] = 0;rain_draw[35][96] = 0;rain_draw[36][96] = 0;rain_draw[37][96] = 0;rain_draw[38][96] = 0;rain_draw[39][96] = 0;rain_draw[40][96] = 0;rain_draw[41][96] = 0;rain_draw[42][96] = 0;rain_draw[43][96] = 0;rain_draw[44][96] = 0;rain_draw[45][96] = 0;rain_draw[46][96] = 0;rain_draw[47][96] = 0;rain_draw[48][96] = 0;rain_draw[49][96] = 0;rain_draw[50][96] = 0;rain_draw[51][96] = 0;rain_draw[52][96] = 0;rain_draw[53][96] = 0;rain_draw[54][96] = 0;rain_draw[55][96] = 0;rain_draw[56][96] = 0;rain_draw[57][96] = 0;rain_draw[58][96] = 0;rain_draw[59][96] = 0;rain_draw[60][96] = 0;rain_draw[61][96] = 0;rain_draw[62][96] = 0;rain_draw[63][96] = 0;rain_draw[64][96] = 0;rain_draw[65][96] = 0;rain_draw[66][96] = 0;rain_draw[67][96] = 0;rain_draw[68][96] = 0;rain_draw[69][96] = 0;rain_draw[70][96] = 0;rain_draw[71][96] = 0;rain_draw[72][96] = 0;rain_draw[73][96] = 0;rain_draw[74][96] = 0;rain_draw[75][96] = 0;rain_draw[76][96] = 0;rain_draw[77][96] = 0;rain_draw[78][96] = 0;rain_draw[79][96] = 0;rain_draw[80][96] = 0;rain_draw[81][96] = 0;rain_draw[82][96] = 0;rain_draw[83][96] = 0;rain_draw[84][96] = 0;rain_draw[85][96] = 0;rain_draw[86][96] = 0;rain_draw[87][96] = 0;rain_draw[88][96] = 0;rain_draw[89][96] = 0;rain_draw[90][96] = 0;rain_draw[91][96] = 0;rain_draw[92][96] = 0;rain_draw[93][96] = 0;rain_draw[94][96] = 0;rain_draw[95][96] = 0;
        rain_draw[0][97] = 0;rain_draw[1][97] = 0;rain_draw[2][97] = 0;rain_draw[3][97] = 0;rain_draw[4][97] = 0;rain_draw[5][97] = 0;rain_draw[6][97] = 1;rain_draw[7][97] = 1;rain_draw[8][97] = 1;rain_draw[9][97] = 0;rain_draw[10][97] = 0;rain_draw[11][97] = 0;rain_draw[12][97] = 0;rain_draw[13][97] = 0;rain_draw[14][97] = 0;rain_draw[15][97] = 0;rain_draw[16][97] = 0;rain_draw[17][97] = 0;rain_draw[18][97] = 0;rain_draw[19][97] = 0;rain_draw[20][97] = 0;rain_draw[21][97] = 0;rain_draw[22][97] = 0;rain_draw[23][97] = 0;rain_draw[24][97] = 0;rain_draw[25][97] = 0;rain_draw[26][97] = 0;rain_draw[27][97] = 0;rain_draw[28][97] = 0;rain_draw[29][97] = 0;rain_draw[30][97] = 0;rain_draw[31][97] = 0;rain_draw[32][97] = 0;rain_draw[33][97] = 0;rain_draw[34][97] = 0;rain_draw[35][97] = 0;rain_draw[36][97] = 0;rain_draw[37][97] = 0;rain_draw[38][97] = 0;rain_draw[39][97] = 0;rain_draw[40][97] = 0;rain_draw[41][97] = 0;rain_draw[42][97] = 0;rain_draw[43][97] = 0;rain_draw[44][97] = 0;rain_draw[45][97] = 0;rain_draw[46][97] = 0;rain_draw[47][97] = 0;rain_draw[48][97] = 0;rain_draw[49][97] = 0;rain_draw[50][97] = 0;rain_draw[51][97] = 0;rain_draw[52][97] = 0;rain_draw[53][97] = 0;rain_draw[54][97] = 0;rain_draw[55][97] = 0;rain_draw[56][97] = 0;rain_draw[57][97] = 0;rain_draw[58][97] = 0;rain_draw[59][97] = 0;rain_draw[60][97] = 0;rain_draw[61][97] = 0;rain_draw[62][97] = 0;rain_draw[63][97] = 0;rain_draw[64][97] = 0;rain_draw[65][97] = 0;rain_draw[66][97] = 0;rain_draw[67][97] = 0;rain_draw[68][97] = 0;rain_draw[69][97] = 0;rain_draw[70][97] = 0;rain_draw[71][97] = 0;rain_draw[72][97] = 0;rain_draw[73][97] = 0;rain_draw[74][97] = 0;rain_draw[75][97] = 0;rain_draw[76][97] = 0;rain_draw[77][97] = 0;rain_draw[78][97] = 0;rain_draw[79][97] = 0;rain_draw[80][97] = 0;rain_draw[81][97] = 0;rain_draw[82][97] = 0;rain_draw[83][97] = 0;rain_draw[84][97] = 0;rain_draw[85][97] = 0;rain_draw[86][97] = 0;rain_draw[87][97] = 0;rain_draw[88][97] = 0;rain_draw[89][97] = 0;rain_draw[90][97] = 0;rain_draw[91][97] = 0;rain_draw[92][97] = 0;rain_draw[93][97] = 0;rain_draw[94][97] = 0;rain_draw[95][97] = 0;
        rain_draw[0][98] = 0;rain_draw[1][98] = 0;rain_draw[2][98] = 0;rain_draw[3][98] = 0;rain_draw[4][98] = 0;rain_draw[5][98] = 1;rain_draw[6][98] = 1;rain_draw[7][98] = 1;rain_draw[8][98] = 0;rain_draw[9][98] = 0;rain_draw[10][98] = 0;rain_draw[11][98] = 0;rain_draw[12][98] = 0;rain_draw[13][98] = 0;rain_draw[14][98] = 0;rain_draw[15][98] = 0;rain_draw[16][98] = 0;rain_draw[17][98] = 0;rain_draw[18][98] = 0;rain_draw[19][98] = 0;rain_draw[20][98] = 0;rain_draw[21][98] = 0;rain_draw[22][98] = 0;rain_draw[23][98] = 0;rain_draw[24][98] = 0;rain_draw[25][98] = 0;rain_draw[26][98] = 0;rain_draw[27][98] = 0;rain_draw[28][98] = 0;rain_draw[29][98] = 0;rain_draw[30][98] = 0;rain_draw[31][98] = 0;rain_draw[32][98] = 0;rain_draw[33][98] = 0;rain_draw[34][98] = 0;rain_draw[35][98] = 0;rain_draw[36][98] = 0;rain_draw[37][98] = 0;rain_draw[38][98] = 0;rain_draw[39][98] = 0;rain_draw[40][98] = 0;rain_draw[41][98] = 0;rain_draw[42][98] = 0;rain_draw[43][98] = 0;rain_draw[44][98] = 0;rain_draw[45][98] = 0;rain_draw[46][98] = 0;rain_draw[47][98] = 0;rain_draw[48][98] = 0;rain_draw[49][98] = 0;rain_draw[50][98] = 0;rain_draw[51][98] = 0;rain_draw[52][98] = 0;rain_draw[53][98] = 0;rain_draw[54][98] = 0;rain_draw[55][98] = 0;rain_draw[56][98] = 0;rain_draw[57][98] = 0;rain_draw[58][98] = 0;rain_draw[59][98] = 0;rain_draw[60][98] = 0;rain_draw[61][98] = 0;rain_draw[62][98] = 0;rain_draw[63][98] = 0;rain_draw[64][98] = 0;rain_draw[65][98] = 0;rain_draw[66][98] = 0;rain_draw[67][98] = 0;rain_draw[68][98] = 0;rain_draw[69][98] = 0;rain_draw[70][98] = 0;rain_draw[71][98] = 0;rain_draw[72][98] = 0;rain_draw[73][98] = 0;rain_draw[74][98] = 0;rain_draw[75][98] = 0;rain_draw[76][98] = 0;rain_draw[77][98] = 0;rain_draw[78][98] = 0;rain_draw[79][98] = 0;rain_draw[80][98] = 0;rain_draw[81][98] = 0;rain_draw[82][98] = 0;rain_draw[83][98] = 0;rain_draw[84][98] = 0;rain_draw[85][98] = 0;rain_draw[86][98] = 0;rain_draw[87][98] = 0;rain_draw[88][98] = 0;rain_draw[89][98] = 0;rain_draw[90][98] = 0;rain_draw[91][98] = 0;rain_draw[92][98] = 0;rain_draw[93][98] = 0;rain_draw[94][98] = 0;rain_draw[95][98] = 0;
        rain_draw[0][99] = 0;rain_draw[1][99] = 0;rain_draw[2][99] = 0;rain_draw[3][99] = 0;rain_draw[4][99] = 1;rain_draw[5][99] = 1;rain_draw[6][99] = 1;rain_draw[7][99] = 0;rain_draw[8][99] = 0;rain_draw[9][99] = 0;rain_draw[10][99] = 0;rain_draw[11][99] = 0;rain_draw[12][99] = 0;rain_draw[13][99] = 0;rain_draw[14][99] = 0;rain_draw[15][99] = 0;rain_draw[16][99] = 0;rain_draw[17][99] = 0;rain_draw[18][99] = 0;rain_draw[19][99] = 0;rain_draw[20][99] = 0;rain_draw[21][99] = 0;rain_draw[22][99] = 0;rain_draw[23][99] = 0;rain_draw[24][99] = 0;rain_draw[25][99] = 0;rain_draw[26][99] = 0;rain_draw[27][99] = 0;rain_draw[28][99] = 0;rain_draw[29][99] = 0;rain_draw[30][99] = 0;rain_draw[31][99] = 0;rain_draw[32][99] = 0;rain_draw[33][99] = 0;rain_draw[34][99] = 0;rain_draw[35][99] = 0;rain_draw[36][99] = 0;rain_draw[37][99] = 0;rain_draw[38][99] = 0;rain_draw[39][99] = 0;rain_draw[40][99] = 0;rain_draw[41][99] = 0;rain_draw[42][99] = 0;rain_draw[43][99] = 0;rain_draw[44][99] = 0;rain_draw[45][99] = 0;rain_draw[46][99] = 0;rain_draw[47][99] = 0;rain_draw[48][99] = 0;rain_draw[49][99] = 0;rain_draw[50][99] = 0;rain_draw[51][99] = 0;rain_draw[52][99] = 0;rain_draw[53][99] = 0;rain_draw[54][99] = 0;rain_draw[55][99] = 0;rain_draw[56][99] = 0;rain_draw[57][99] = 0;rain_draw[58][99] = 0;rain_draw[59][99] = 0;rain_draw[60][99] = 0;rain_draw[61][99] = 0;rain_draw[62][99] = 0;rain_draw[63][99] = 0;rain_draw[64][99] = 0;rain_draw[65][99] = 0;rain_draw[66][99] = 0;rain_draw[67][99] = 0;rain_draw[68][99] = 0;rain_draw[69][99] = 0;rain_draw[70][99] = 0;rain_draw[71][99] = 0;rain_draw[72][99] = 0;rain_draw[73][99] = 0;rain_draw[74][99] = 0;rain_draw[75][99] = 0;rain_draw[76][99] = 0;rain_draw[77][99] = 0;rain_draw[78][99] = 0;rain_draw[79][99] = 0;rain_draw[80][99] = 0;rain_draw[81][99] = 0;rain_draw[82][99] = 0;rain_draw[83][99] = 0;rain_draw[84][99] = 0;rain_draw[85][99] = 0;rain_draw[86][99] = 0;rain_draw[87][99] = 0;rain_draw[88][99] = 0;rain_draw[89][99] = 0;rain_draw[90][99] = 0;rain_draw[91][99] = 0;rain_draw[92][99] = 0;rain_draw[93][99] = 0;rain_draw[94][99] = 0;rain_draw[95][99] = 0;
        rain_draw[0][100] = 0;rain_draw[1][100] = 0;rain_draw[2][100] = 0;rain_draw[3][100] = 1;rain_draw[4][100] = 1;rain_draw[5][100] = 1;rain_draw[6][100] = 0;rain_draw[7][100] = 0;rain_draw[8][100] = 0;rain_draw[9][100] = 0;rain_draw[10][100] = 0;rain_draw[11][100] = 0;rain_draw[12][100] = 0;rain_draw[13][100] = 0;rain_draw[14][100] = 0;rain_draw[15][100] = 0;rain_draw[16][100] = 0;rain_draw[17][100] = 0;rain_draw[18][100] = 0;rain_draw[19][100] = 0;rain_draw[20][100] = 0;rain_draw[21][100] = 0;rain_draw[22][100] = 0;rain_draw[23][100] = 0;rain_draw[24][100] = 0;rain_draw[25][100] = 0;rain_draw[26][100] = 0;rain_draw[27][100] = 0;rain_draw[28][100] = 0;rain_draw[29][100] = 0;rain_draw[30][100] = 0;rain_draw[31][100] = 0;rain_draw[32][100] = 0;rain_draw[33][100] = 0;rain_draw[34][100] = 0;rain_draw[35][100] = 0;rain_draw[36][100] = 0;rain_draw[37][100] = 0;rain_draw[38][100] = 0;rain_draw[39][100] = 0;rain_draw[40][100] = 0;rain_draw[41][100] = 0;rain_draw[42][100] = 0;rain_draw[43][100] = 0;rain_draw[44][100] = 0;rain_draw[45][100] = 0;rain_draw[46][100] = 0;rain_draw[47][100] = 0;rain_draw[48][100] = 0;rain_draw[49][100] = 0;rain_draw[50][100] = 0;rain_draw[51][100] = 0;rain_draw[52][100] = 0;rain_draw[53][100] = 0;rain_draw[54][100] = 0;rain_draw[55][100] = 0;rain_draw[56][100] = 0;rain_draw[57][100] = 0;rain_draw[58][100] = 0;rain_draw[59][100] = 0;rain_draw[60][100] = 0;rain_draw[61][100] = 0;rain_draw[62][100] = 0;rain_draw[63][100] = 0;rain_draw[64][100] = 0;rain_draw[65][100] = 0;rain_draw[66][100] = 0;rain_draw[67][100] = 0;rain_draw[68][100] = 0;rain_draw[69][100] = 0;rain_draw[70][100] = 0;rain_draw[71][100] = 0;rain_draw[72][100] = 0;rain_draw[73][100] = 0;rain_draw[74][100] = 0;rain_draw[75][100] = 0;rain_draw[76][100] = 0;rain_draw[77][100] = 0;rain_draw[78][100] = 0;rain_draw[79][100] = 0;rain_draw[80][100] = 0;rain_draw[81][100] = 0;rain_draw[82][100] = 0;rain_draw[83][100] = 0;rain_draw[84][100] = 0;rain_draw[85][100] = 0;rain_draw[86][100] = 0;rain_draw[87][100] = 0;rain_draw[88][100] = 0;rain_draw[89][100] = 0;rain_draw[90][100] = 0;rain_draw[91][100] = 0;rain_draw[92][100] = 0;rain_draw[93][100] = 0;rain_draw[94][100] = 0;rain_draw[95][100] = 0;
        rain_draw[0][101] = 0;rain_draw[1][101] = 0;rain_draw[2][101] = 0;rain_draw[3][101] = 0;rain_draw[4][101] = 0;rain_draw[5][101] = 0;rain_draw[6][101] = 0;rain_draw[7][101] = 0;rain_draw[8][101] = 0;rain_draw[9][101] = 0;rain_draw[10][101] = 0;rain_draw[11][101] = 0;rain_draw[12][101] = 0;rain_draw[13][101] = 0;rain_draw[14][101] = 0;rain_draw[15][101] = 0;rain_draw[16][101] = 0;rain_draw[17][101] = 0;rain_draw[18][101] = 0;rain_draw[19][101] = 0;rain_draw[20][101] = 0;rain_draw[21][101] = 0;rain_draw[22][101] = 0;rain_draw[23][101] = 0;rain_draw[24][101] = 0;rain_draw[25][101] = 0;rain_draw[26][101] = 0;rain_draw[27][101] = 0;rain_draw[28][101] = 0;rain_draw[29][101] = 0;rain_draw[30][101] = 0;rain_draw[31][101] = 0;rain_draw[32][101] = 0;rain_draw[33][101] = 0;rain_draw[34][101] = 0;rain_draw[35][101] = 0;rain_draw[36][101] = 0;rain_draw[37][101] = 0;rain_draw[38][101] = 0;rain_draw[39][101] = 0;rain_draw[40][101] = 0;rain_draw[41][101] = 0;rain_draw[42][101] = 0;rain_draw[43][101] = 0;rain_draw[44][101] = 0;rain_draw[45][101] = 0;rain_draw[46][101] = 0;rain_draw[47][101] = 0;rain_draw[48][101] = 0;rain_draw[49][101] = 0;rain_draw[50][101] = 0;rain_draw[51][101] = 0;rain_draw[52][101] = 0;rain_draw[53][101] = 0;rain_draw[54][101] = 0;rain_draw[55][101] = 0;rain_draw[56][101] = 0;rain_draw[57][101] = 0;rain_draw[58][101] = 0;rain_draw[59][101] = 0;rain_draw[60][101] = 0;rain_draw[61][101] = 0;rain_draw[62][101] = 0;rain_draw[63][101] = 0;rain_draw[64][101] = 0;rain_draw[65][101] = 0;rain_draw[66][101] = 0;rain_draw[67][101] = 0;rain_draw[68][101] = 0;rain_draw[69][101] = 0;rain_draw[70][101] = 0;rain_draw[71][101] = 0;rain_draw[72][101] = 0;rain_draw[73][101] = 0;rain_draw[74][101] = 0;rain_draw[75][101] = 0;rain_draw[76][101] = 0;rain_draw[77][101] = 0;rain_draw[78][101] = 0;rain_draw[79][101] = 0;rain_draw[80][101] = 0;rain_draw[81][101] = 0;rain_draw[82][101] = 0;rain_draw[83][101] = 0;rain_draw[84][101] = 0;rain_draw[85][101] = 0;rain_draw[86][101] = 0;rain_draw[87][101] = 0;rain_draw[88][101] = 0;rain_draw[89][101] = 0;rain_draw[90][101] = 0;rain_draw[91][101] = 0;rain_draw[92][101] = 0;rain_draw[93][101] = 0;rain_draw[94][101] = 0;rain_draw[95][101] = 0;
        rain_draw[0][102] = 0;rain_draw[1][102] = 0;rain_draw[2][102] = 0;rain_draw[3][102] = 0;rain_draw[4][102] = 0;rain_draw[5][102] = 0;rain_draw[6][102] = 0;rain_draw[7][102] = 0;rain_draw[8][102] = 0;rain_draw[9][102] = 0;rain_draw[10][102] = 0;rain_draw[11][102] = 0;rain_draw[12][102] = 0;rain_draw[13][102] = 0;rain_draw[14][102] = 0;rain_draw[15][102] = 0;rain_draw[16][102] = 0;rain_draw[17][102] = 0;rain_draw[18][102] = 0;rain_draw[19][102] = 0;rain_draw[20][102] = 0;rain_draw[21][102] = 0;rain_draw[22][102] = 0;rain_draw[23][102] = 0;rain_draw[24][102] = 0;rain_draw[25][102] = 0;rain_draw[26][102] = 0;rain_draw[27][102] = 0;rain_draw[28][102] = 0;rain_draw[29][102] = 0;rain_draw[30][102] = 0;rain_draw[31][102] = 0;rain_draw[32][102] = 0;rain_draw[33][102] = 0;rain_draw[34][102] = 0;rain_draw[35][102] = 0;rain_draw[36][102] = 0;rain_draw[37][102] = 0;rain_draw[38][102] = 0;rain_draw[39][102] = 0;rain_draw[40][102] = 0;rain_draw[41][102] = 0;rain_draw[42][102] = 0;rain_draw[43][102] = 0;rain_draw[44][102] = 0;rain_draw[45][102] = 0;rain_draw[46][102] = 0;rain_draw[47][102] = 0;rain_draw[48][102] = 0;rain_draw[49][102] = 0;rain_draw[50][102] = 0;rain_draw[51][102] = 0;rain_draw[52][102] = 0;rain_draw[53][102] = 0;rain_draw[54][102] = 0;rain_draw[55][102] = 0;rain_draw[56][102] = 0;rain_draw[57][102] = 0;rain_draw[58][102] = 0;rain_draw[59][102] = 0;rain_draw[60][102] = 0;rain_draw[61][102] = 0;rain_draw[62][102] = 0;rain_draw[63][102] = 0;rain_draw[64][102] = 0;rain_draw[65][102] = 0;rain_draw[66][102] = 0;rain_draw[67][102] = 0;rain_draw[68][102] = 0;rain_draw[69][102] = 0;rain_draw[70][102] = 0;rain_draw[71][102] = 0;rain_draw[72][102] = 0;rain_draw[73][102] = 0;rain_draw[74][102] = 0;rain_draw[75][102] = 0;rain_draw[76][102] = 0;rain_draw[77][102] = 0;rain_draw[78][102] = 0;rain_draw[79][102] = 0;rain_draw[80][102] = 0;rain_draw[81][102] = 0;rain_draw[82][102] = 0;rain_draw[83][102] = 0;rain_draw[84][102] = 0;rain_draw[85][102] = 0;rain_draw[86][102] = 0;rain_draw[87][102] = 0;rain_draw[88][102] = 0;rain_draw[89][102] = 0;rain_draw[90][102] = 0;rain_draw[91][102] = 0;rain_draw[92][102] = 0;rain_draw[93][102] = 0;rain_draw[94][102] = 0;rain_draw[95][102] = 0;
        rain_draw[0][103] = 0;rain_draw[1][103] = 0;rain_draw[2][103] = 0;rain_draw[3][103] = 0;rain_draw[4][103] = 0;rain_draw[5][103] = 0;rain_draw[6][103] = 0;rain_draw[7][103] = 0;rain_draw[8][103] = 0;rain_draw[9][103] = 0;rain_draw[10][103] = 0;rain_draw[11][103] = 0;rain_draw[12][103] = 0;rain_draw[13][103] = 0;rain_draw[14][103] = 0;rain_draw[15][103] = 0;rain_draw[16][103] = 0;rain_draw[17][103] = 0;rain_draw[18][103] = 0;rain_draw[19][103] = 0;rain_draw[20][103] = 0;rain_draw[21][103] = 0;rain_draw[22][103] = 0;rain_draw[23][103] = 0;rain_draw[24][103] = 0;rain_draw[25][103] = 0;rain_draw[26][103] = 0;rain_draw[27][103] = 0;rain_draw[28][103] = 0;rain_draw[29][103] = 0;rain_draw[30][103] = 0;rain_draw[31][103] = 0;rain_draw[32][103] = 0;rain_draw[33][103] = 0;rain_draw[34][103] = 0;rain_draw[35][103] = 0;rain_draw[36][103] = 0;rain_draw[37][103] = 0;rain_draw[38][103] = 0;rain_draw[39][103] = 0;rain_draw[40][103] = 0;rain_draw[41][103] = 0;rain_draw[42][103] = 0;rain_draw[43][103] = 0;rain_draw[44][103] = 0;rain_draw[45][103] = 0;rain_draw[46][103] = 0;rain_draw[47][103] = 0;rain_draw[48][103] = 0;rain_draw[49][103] = 0;rain_draw[50][103] = 0;rain_draw[51][103] = 0;rain_draw[52][103] = 0;rain_draw[53][103] = 0;rain_draw[54][103] = 0;rain_draw[55][103] = 0;rain_draw[56][103] = 0;rain_draw[57][103] = 0;rain_draw[58][103] = 0;rain_draw[59][103] = 0;rain_draw[60][103] = 0;rain_draw[61][103] = 0;rain_draw[62][103] = 0;rain_draw[63][103] = 0;rain_draw[64][103] = 0;rain_draw[65][103] = 0;rain_draw[66][103] = 0;rain_draw[67][103] = 0;rain_draw[68][103] = 0;rain_draw[69][103] = 0;rain_draw[70][103] = 0;rain_draw[71][103] = 0;rain_draw[72][103] = 0;rain_draw[73][103] = 0;rain_draw[74][103] = 0;rain_draw[75][103] = 0;rain_draw[76][103] = 0;rain_draw[77][103] = 0;rain_draw[78][103] = 0;rain_draw[79][103] = 0;rain_draw[80][103] = 0;rain_draw[81][103] = 0;rain_draw[82][103] = 0;rain_draw[83][103] = 0;rain_draw[84][103] = 0;rain_draw[85][103] = 0;rain_draw[86][103] = 0;rain_draw[87][103] = 0;rain_draw[88][103] = 0;rain_draw[89][103] = 0;rain_draw[90][103] = 0;rain_draw[91][103] = 0;rain_draw[92][103] = 0;rain_draw[93][103] = 0;rain_draw[94][103] = 0;rain_draw[95][103] = 0;
        rain_draw[0][104] = 0;rain_draw[1][104] = 0;rain_draw[2][104] = 0;rain_draw[3][104] = 0;rain_draw[4][104] = 0;rain_draw[5][104] = 0;rain_draw[6][104] = 0;rain_draw[7][104] = 0;rain_draw[8][104] = 0;rain_draw[9][104] = 0;rain_draw[10][104] = 0;rain_draw[11][104] = 0;rain_draw[12][104] = 0;rain_draw[13][104] = 0;rain_draw[14][104] = 0;rain_draw[15][104] = 0;rain_draw[16][104] = 0;rain_draw[17][104] = 0;rain_draw[18][104] = 0;rain_draw[19][104] = 0;rain_draw[20][104] = 0;rain_draw[21][104] = 0;rain_draw[22][104] = 0;rain_draw[23][104] = 0;rain_draw[24][104] = 0;rain_draw[25][104] = 0;rain_draw[26][104] = 0;rain_draw[27][104] = 0;rain_draw[28][104] = 0;rain_draw[29][104] = 0;rain_draw[30][104] = 0;rain_draw[31][104] = 0;rain_draw[32][104] = 0;rain_draw[33][104] = 0;rain_draw[34][104] = 0;rain_draw[35][104] = 0;rain_draw[36][104] = 0;rain_draw[37][104] = 0;rain_draw[38][104] = 0;rain_draw[39][104] = 0;rain_draw[40][104] = 0;rain_draw[41][104] = 0;rain_draw[42][104] = 0;rain_draw[43][104] = 0;rain_draw[44][104] = 0;rain_draw[45][104] = 0;rain_draw[46][104] = 0;rain_draw[47][104] = 0;rain_draw[48][104] = 0;rain_draw[49][104] = 0;rain_draw[50][104] = 0;rain_draw[51][104] = 0;rain_draw[52][104] = 0;rain_draw[53][104] = 0;rain_draw[54][104] = 0;rain_draw[55][104] = 0;rain_draw[56][104] = 0;rain_draw[57][104] = 0;rain_draw[58][104] = 0;rain_draw[59][104] = 0;rain_draw[60][104] = 0;rain_draw[61][104] = 0;rain_draw[62][104] = 0;rain_draw[63][104] = 0;rain_draw[64][104] = 0;rain_draw[65][104] = 0;rain_draw[66][104] = 0;rain_draw[67][104] = 0;rain_draw[68][104] = 0;rain_draw[69][104] = 0;rain_draw[70][104] = 0;rain_draw[71][104] = 0;rain_draw[72][104] = 0;rain_draw[73][104] = 0;rain_draw[74][104] = 0;rain_draw[75][104] = 0;rain_draw[76][104] = 0;rain_draw[77][104] = 0;rain_draw[78][104] = 0;rain_draw[79][104] = 0;rain_draw[80][104] = 0;rain_draw[81][104] = 0;rain_draw[82][104] = 0;rain_draw[83][104] = 0;rain_draw[84][104] = 0;rain_draw[85][104] = 0;rain_draw[86][104] = 0;rain_draw[87][104] = 0;rain_draw[88][104] = 0;rain_draw[89][104] = 0;rain_draw[90][104] = 0;rain_draw[91][104] = 0;rain_draw[92][104] = 0;rain_draw[93][104] = 0;rain_draw[94][104] = 0;rain_draw[95][104] = 0;
        rain_draw[0][105] = 0;rain_draw[1][105] = 0;rain_draw[2][105] = 0;rain_draw[3][105] = 0;rain_draw[4][105] = 0;rain_draw[5][105] = 0;rain_draw[6][105] = 0;rain_draw[7][105] = 0;rain_draw[8][105] = 0;rain_draw[9][105] = 0;rain_draw[10][105] = 0;rain_draw[11][105] = 0;rain_draw[12][105] = 0;rain_draw[13][105] = 0;rain_draw[14][105] = 0;rain_draw[15][105] = 0;rain_draw[16][105] = 0;rain_draw[17][105] = 0;rain_draw[18][105] = 0;rain_draw[19][105] = 0;rain_draw[20][105] = 0;rain_draw[21][105] = 0;rain_draw[22][105] = 0;rain_draw[23][105] = 0;rain_draw[24][105] = 0;rain_draw[25][105] = 0;rain_draw[26][105] = 0;rain_draw[27][105] = 0;rain_draw[28][105] = 0;rain_draw[29][105] = 0;rain_draw[30][105] = 0;rain_draw[31][105] = 0;rain_draw[32][105] = 0;rain_draw[33][105] = 0;rain_draw[34][105] = 0;rain_draw[35][105] = 0;rain_draw[36][105] = 0;rain_draw[37][105] = 0;rain_draw[38][105] = 0;rain_draw[39][105] = 0;rain_draw[40][105] = 0;rain_draw[41][105] = 0;rain_draw[42][105] = 0;rain_draw[43][105] = 0;rain_draw[44][105] = 0;rain_draw[45][105] = 0;rain_draw[46][105] = 0;rain_draw[47][105] = 0;rain_draw[48][105] = 0;rain_draw[49][105] = 0;rain_draw[50][105] = 0;rain_draw[51][105] = 0;rain_draw[52][105] = 0;rain_draw[53][105] = 0;rain_draw[54][105] = 0;rain_draw[55][105] = 0;rain_draw[56][105] = 0;rain_draw[57][105] = 0;rain_draw[58][105] = 0;rain_draw[59][105] = 0;rain_draw[60][105] = 0;rain_draw[61][105] = 0;rain_draw[62][105] = 0;rain_draw[63][105] = 0;rain_draw[64][105] = 0;rain_draw[65][105] = 0;rain_draw[66][105] = 0;rain_draw[67][105] = 1;rain_draw[68][105] = 1;rain_draw[69][105] = 1;rain_draw[70][105] = 0;rain_draw[71][105] = 0;rain_draw[72][105] = 0;rain_draw[73][105] = 0;rain_draw[74][105] = 0;rain_draw[75][105] = 0;rain_draw[76][105] = 0;rain_draw[77][105] = 0;rain_draw[78][105] = 0;rain_draw[79][105] = 0;rain_draw[80][105] = 0;rain_draw[81][105] = 0;rain_draw[82][105] = 0;rain_draw[83][105] = 0;rain_draw[84][105] = 0;rain_draw[85][105] = 0;rain_draw[86][105] = 0;rain_draw[87][105] = 0;rain_draw[88][105] = 0;rain_draw[89][105] = 0;rain_draw[90][105] = 0;rain_draw[91][105] = 0;rain_draw[92][105] = 0;rain_draw[93][105] = 0;rain_draw[94][105] = 0;rain_draw[95][105] = 0;
        rain_draw[0][106] = 0;rain_draw[1][106] = 0;rain_draw[2][106] = 0;rain_draw[3][106] = 0;rain_draw[4][106] = 0;rain_draw[5][106] = 0;rain_draw[6][106] = 0;rain_draw[7][106] = 0;rain_draw[8][106] = 0;rain_draw[9][106] = 0;rain_draw[10][106] = 0;rain_draw[11][106] = 0;rain_draw[12][106] = 0;rain_draw[13][106] = 0;rain_draw[14][106] = 0;rain_draw[15][106] = 0;rain_draw[16][106] = 0;rain_draw[17][106] = 0;rain_draw[18][106] = 0;rain_draw[19][106] = 0;rain_draw[20][106] = 0;rain_draw[21][106] = 0;rain_draw[22][106] = 0;rain_draw[23][106] = 0;rain_draw[24][106] = 0;rain_draw[25][106] = 0;rain_draw[26][106] = 0;rain_draw[27][106] = 0;rain_draw[28][106] = 0;rain_draw[29][106] = 0;rain_draw[30][106] = 0;rain_draw[31][106] = 0;rain_draw[32][106] = 0;rain_draw[33][106] = 0;rain_draw[34][106] = 0;rain_draw[35][106] = 0;rain_draw[36][106] = 0;rain_draw[37][106] = 0;rain_draw[38][106] = 0;rain_draw[39][106] = 0;rain_draw[40][106] = 0;rain_draw[41][106] = 0;rain_draw[42][106] = 0;rain_draw[43][106] = 0;rain_draw[44][106] = 0;rain_draw[45][106] = 0;rain_draw[46][106] = 0;rain_draw[47][106] = 0;rain_draw[48][106] = 0;rain_draw[49][106] = 0;rain_draw[50][106] = 0;rain_draw[51][106] = 0;rain_draw[52][106] = 0;rain_draw[53][106] = 0;rain_draw[54][106] = 0;rain_draw[55][106] = 0;rain_draw[56][106] = 0;rain_draw[57][106] = 0;rain_draw[58][106] = 0;rain_draw[59][106] = 0;rain_draw[60][106] = 0;rain_draw[61][106] = 0;rain_draw[62][106] = 0;rain_draw[63][106] = 0;rain_draw[64][106] = 0;rain_draw[65][106] = 0;rain_draw[66][106] = 1;rain_draw[67][106] = 1;rain_draw[68][106] = 1;rain_draw[69][106] = 0;rain_draw[70][106] = 0;rain_draw[71][106] = 0;rain_draw[72][106] = 0;rain_draw[73][106] = 0;rain_draw[74][106] = 0;rain_draw[75][106] = 0;rain_draw[76][106] = 0;rain_draw[77][106] = 0;rain_draw[78][106] = 0;rain_draw[79][106] = 0;rain_draw[80][106] = 0;rain_draw[81][106] = 0;rain_draw[82][106] = 0;rain_draw[83][106] = 0;rain_draw[84][106] = 0;rain_draw[85][106] = 0;rain_draw[86][106] = 0;rain_draw[87][106] = 0;rain_draw[88][106] = 0;rain_draw[89][106] = 0;rain_draw[90][106] = 0;rain_draw[91][106] = 0;rain_draw[92][106] = 0;rain_draw[93][106] = 0;rain_draw[94][106] = 0;rain_draw[95][106] = 0;
        rain_draw[0][107] = 0;rain_draw[1][107] = 0;rain_draw[2][107] = 0;rain_draw[3][107] = 0;rain_draw[4][107] = 0;rain_draw[5][107] = 0;rain_draw[6][107] = 0;rain_draw[7][107] = 0;rain_draw[8][107] = 0;rain_draw[9][107] = 0;rain_draw[10][107] = 0;rain_draw[11][107] = 0;rain_draw[12][107] = 0;rain_draw[13][107] = 0;rain_draw[14][107] = 0;rain_draw[15][107] = 0;rain_draw[16][107] = 0;rain_draw[17][107] = 0;rain_draw[18][107] = 0;rain_draw[19][107] = 0;rain_draw[20][107] = 0;rain_draw[21][107] = 0;rain_draw[22][107] = 0;rain_draw[23][107] = 0;rain_draw[24][107] = 0;rain_draw[25][107] = 0;rain_draw[26][107] = 0;rain_draw[27][107] = 0;rain_draw[28][107] = 0;rain_draw[29][107] = 0;rain_draw[30][107] = 0;rain_draw[31][107] = 0;rain_draw[32][107] = 0;rain_draw[33][107] = 0;rain_draw[34][107] = 0;rain_draw[35][107] = 0;rain_draw[36][107] = 0;rain_draw[37][107] = 0;rain_draw[38][107] = 0;rain_draw[39][107] = 0;rain_draw[40][107] = 0;rain_draw[41][107] = 0;rain_draw[42][107] = 0;rain_draw[43][107] = 0;rain_draw[44][107] = 0;rain_draw[45][107] = 0;rain_draw[46][107] = 0;rain_draw[47][107] = 0;rain_draw[48][107] = 0;rain_draw[49][107] = 0;rain_draw[50][107] = 0;rain_draw[51][107] = 0;rain_draw[52][107] = 0;rain_draw[53][107] = 0;rain_draw[54][107] = 0;rain_draw[55][107] = 0;rain_draw[56][107] = 0;rain_draw[57][107] = 0;rain_draw[58][107] = 0;rain_draw[59][107] = 0;rain_draw[60][107] = 0;rain_draw[61][107] = 0;rain_draw[62][107] = 0;rain_draw[63][107] = 0;rain_draw[64][107] = 0;rain_draw[65][107] = 1;rain_draw[66][107] = 1;rain_draw[67][107] = 1;rain_draw[68][107] = 0;rain_draw[69][107] = 0;rain_draw[70][107] = 0;rain_draw[71][107] = 0;rain_draw[72][107] = 0;rain_draw[73][107] = 0;rain_draw[74][107] = 0;rain_draw[75][107] = 0;rain_draw[76][107] = 0;rain_draw[77][107] = 0;rain_draw[78][107] = 0;rain_draw[79][107] = 0;rain_draw[80][107] = 0;rain_draw[81][107] = 0;rain_draw[82][107] = 0;rain_draw[83][107] = 0;rain_draw[84][107] = 0;rain_draw[85][107] = 0;rain_draw[86][107] = 1;rain_draw[87][107] = 1;rain_draw[88][107] = 1;rain_draw[89][107] = 0;rain_draw[90][107] = 0;rain_draw[91][107] = 0;rain_draw[92][107] = 0;rain_draw[93][107] = 0;rain_draw[94][107] = 0;rain_draw[95][107] = 0;
        rain_draw[0][108] = 0;rain_draw[1][108] = 0;rain_draw[2][108] = 0;rain_draw[3][108] = 0;rain_draw[4][108] = 0;rain_draw[5][108] = 0;rain_draw[6][108] = 0;rain_draw[7][108] = 0;rain_draw[8][108] = 0;rain_draw[9][108] = 0;rain_draw[10][108] = 0;rain_draw[11][108] = 0;rain_draw[12][108] = 0;rain_draw[13][108] = 0;rain_draw[14][108] = 0;rain_draw[15][108] = 0;rain_draw[16][108] = 0;rain_draw[17][108] = 0;rain_draw[18][108] = 0;rain_draw[19][108] = 0;rain_draw[20][108] = 0;rain_draw[21][108] = 0;rain_draw[22][108] = 0;rain_draw[23][108] = 0;rain_draw[24][108] = 0;rain_draw[25][108] = 0;rain_draw[26][108] = 0;rain_draw[27][108] = 1;rain_draw[28][108] = 1;rain_draw[29][108] = 1;rain_draw[30][108] = 0;rain_draw[31][108] = 0;rain_draw[32][108] = 0;rain_draw[33][108] = 0;rain_draw[34][108] = 0;rain_draw[35][108] = 0;rain_draw[36][108] = 0;rain_draw[37][108] = 0;rain_draw[38][108] = 0;rain_draw[39][108] = 0;rain_draw[40][108] = 0;rain_draw[41][108] = 0;rain_draw[42][108] = 0;rain_draw[43][108] = 0;rain_draw[44][108] = 0;rain_draw[45][108] = 0;rain_draw[46][108] = 0;rain_draw[47][108] = 0;rain_draw[48][108] = 0;rain_draw[49][108] = 0;rain_draw[50][108] = 0;rain_draw[51][108] = 0;rain_draw[52][108] = 0;rain_draw[53][108] = 0;rain_draw[54][108] = 0;rain_draw[55][108] = 0;rain_draw[56][108] = 0;rain_draw[57][108] = 0;rain_draw[58][108] = 0;rain_draw[59][108] = 0;rain_draw[60][108] = 0;rain_draw[61][108] = 0;rain_draw[62][108] = 0;rain_draw[63][108] = 0;rain_draw[64][108] = 1;rain_draw[65][108] = 1;rain_draw[66][108] = 1;rain_draw[67][108] = 0;rain_draw[68][108] = 0;rain_draw[69][108] = 0;rain_draw[70][108] = 0;rain_draw[71][108] = 0;rain_draw[72][108] = 0;rain_draw[73][108] = 0;rain_draw[74][108] = 0;rain_draw[75][108] = 0;rain_draw[76][108] = 0;rain_draw[77][108] = 0;rain_draw[78][108] = 0;rain_draw[79][108] = 0;rain_draw[80][108] = 0;rain_draw[81][108] = 0;rain_draw[82][108] = 0;rain_draw[83][108] = 0;rain_draw[84][108] = 0;rain_draw[85][108] = 1;rain_draw[86][108] = 1;rain_draw[87][108] = 1;rain_draw[88][108] = 0;rain_draw[89][108] = 0;rain_draw[90][108] = 0;rain_draw[91][108] = 0;rain_draw[92][108] = 0;rain_draw[93][108] = 0;rain_draw[94][108] = 0;rain_draw[95][108] = 0;
        rain_draw[0][109] = 0;rain_draw[1][109] = 0;rain_draw[2][109] = 0;rain_draw[3][109] = 0;rain_draw[4][109] = 0;rain_draw[5][109] = 0;rain_draw[6][109] = 0;rain_draw[7][109] = 0;rain_draw[8][109] = 0;rain_draw[9][109] = 0;rain_draw[10][109] = 0;rain_draw[11][109] = 0;rain_draw[12][109] = 0;rain_draw[13][109] = 0;rain_draw[14][109] = 0;rain_draw[15][109] = 0;rain_draw[16][109] = 0;rain_draw[17][109] = 0;rain_draw[18][109] = 0;rain_draw[19][109] = 0;rain_draw[20][109] = 0;rain_draw[21][109] = 0;rain_draw[22][109] = 0;rain_draw[23][109] = 0;rain_draw[24][109] = 0;rain_draw[25][109] = 0;rain_draw[26][109] = 1;rain_draw[27][109] = 1;rain_draw[28][109] = 1;rain_draw[29][109] = 0;rain_draw[30][109] = 0;rain_draw[31][109] = 0;rain_draw[32][109] = 0;rain_draw[33][109] = 0;rain_draw[34][109] = 0;rain_draw[35][109] = 0;rain_draw[36][109] = 0;rain_draw[37][109] = 0;rain_draw[38][109] = 0;rain_draw[39][109] = 0;rain_draw[40][109] = 0;rain_draw[41][109] = 0;rain_draw[42][109] = 0;rain_draw[43][109] = 0;rain_draw[44][109] = 0;rain_draw[45][109] = 0;rain_draw[46][109] = 0;rain_draw[47][109] = 0;rain_draw[48][109] = 0;rain_draw[49][109] = 0;rain_draw[50][109] = 0;rain_draw[51][109] = 0;rain_draw[52][109] = 0;rain_draw[53][109] = 0;rain_draw[54][109] = 0;rain_draw[55][109] = 0;rain_draw[56][109] = 0;rain_draw[57][109] = 0;rain_draw[58][109] = 0;rain_draw[59][109] = 0;rain_draw[60][109] = 0;rain_draw[61][109] = 0;rain_draw[62][109] = 0;rain_draw[63][109] = 1;rain_draw[64][109] = 1;rain_draw[65][109] = 1;rain_draw[66][109] = 0;rain_draw[67][109] = 0;rain_draw[68][109] = 0;rain_draw[69][109] = 0;rain_draw[70][109] = 0;rain_draw[71][109] = 0;rain_draw[72][109] = 0;rain_draw[73][109] = 0;rain_draw[74][109] = 0;rain_draw[75][109] = 0;rain_draw[76][109] = 0;rain_draw[77][109] = 0;rain_draw[78][109] = 0;rain_draw[79][109] = 0;rain_draw[80][109] = 0;rain_draw[81][109] = 0;rain_draw[82][109] = 0;rain_draw[83][109] = 0;rain_draw[84][109] = 1;rain_draw[85][109] = 1;rain_draw[86][109] = 1;rain_draw[87][109] = 0;rain_draw[88][109] = 0;rain_draw[89][109] = 0;rain_draw[90][109] = 0;rain_draw[91][109] = 0;rain_draw[92][109] = 0;rain_draw[93][109] = 0;rain_draw[94][109] = 0;rain_draw[95][109] = 0;
        rain_draw[0][110] = 0;rain_draw[1][110] = 0;rain_draw[2][110] = 0;rain_draw[3][110] = 0;rain_draw[4][110] = 0;rain_draw[5][110] = 0;rain_draw[6][110] = 0;rain_draw[7][110] = 0;rain_draw[8][110] = 0;rain_draw[9][110] = 0;rain_draw[10][110] = 0;rain_draw[11][110] = 0;rain_draw[12][110] = 0;rain_draw[13][110] = 0;rain_draw[14][110] = 0;rain_draw[15][110] = 0;rain_draw[16][110] = 0;rain_draw[17][110] = 0;rain_draw[18][110] = 0;rain_draw[19][110] = 0;rain_draw[20][110] = 0;rain_draw[21][110] = 0;rain_draw[22][110] = 0;rain_draw[23][110] = 0;rain_draw[24][110] = 0;rain_draw[25][110] = 1;rain_draw[26][110] = 1;rain_draw[27][110] = 1;rain_draw[28][110] = 0;rain_draw[29][110] = 0;rain_draw[30][110] = 0;rain_draw[31][110] = 0;rain_draw[32][110] = 0;rain_draw[33][110] = 0;rain_draw[34][110] = 0;rain_draw[35][110] = 0;rain_draw[36][110] = 0;rain_draw[37][110] = 0;rain_draw[38][110] = 0;rain_draw[39][110] = 0;rain_draw[40][110] = 0;rain_draw[41][110] = 0;rain_draw[42][110] = 0;rain_draw[43][110] = 0;rain_draw[44][110] = 0;rain_draw[45][110] = 0;rain_draw[46][110] = 0;rain_draw[47][110] = 0;rain_draw[48][110] = 0;rain_draw[49][110] = 0;rain_draw[50][110] = 0;rain_draw[51][110] = 0;rain_draw[52][110] = 0;rain_draw[53][110] = 0;rain_draw[54][110] = 0;rain_draw[55][110] = 0;rain_draw[56][110] = 0;rain_draw[57][110] = 0;rain_draw[58][110] = 0;rain_draw[59][110] = 0;rain_draw[60][110] = 0;rain_draw[61][110] = 0;rain_draw[62][110] = 1;rain_draw[63][110] = 1;rain_draw[64][110] = 1;rain_draw[65][110] = 0;rain_draw[66][110] = 0;rain_draw[67][110] = 0;rain_draw[68][110] = 0;rain_draw[69][110] = 0;rain_draw[70][110] = 0;rain_draw[71][110] = 0;rain_draw[72][110] = 0;rain_draw[73][110] = 0;rain_draw[74][110] = 0;rain_draw[75][110] = 0;rain_draw[76][110] = 0;rain_draw[77][110] = 0;rain_draw[78][110] = 0;rain_draw[79][110] = 0;rain_draw[80][110] = 0;rain_draw[81][110] = 0;rain_draw[82][110] = 0;rain_draw[83][110] = 1;rain_draw[84][110] = 1;rain_draw[85][110] = 1;rain_draw[86][110] = 0;rain_draw[87][110] = 0;rain_draw[88][110] = 0;rain_draw[89][110] = 0;rain_draw[90][110] = 0;rain_draw[91][110] = 0;rain_draw[92][110] = 0;rain_draw[93][110] = 0;rain_draw[94][110] = 0;rain_draw[95][110] = 0;
        rain_draw[0][111] = 0;rain_draw[1][111] = 0;rain_draw[2][111] = 0;rain_draw[3][111] = 0;rain_draw[4][111] = 0;rain_draw[5][111] = 0;rain_draw[6][111] = 0;rain_draw[7][111] = 0;rain_draw[8][111] = 0;rain_draw[9][111] = 0;rain_draw[10][111] = 0;rain_draw[11][111] = 0;rain_draw[12][111] = 0;rain_draw[13][111] = 0;rain_draw[14][111] = 0;rain_draw[15][111] = 0;rain_draw[16][111] = 0;rain_draw[17][111] = 0;rain_draw[18][111] = 0;rain_draw[19][111] = 0;rain_draw[20][111] = 0;rain_draw[21][111] = 0;rain_draw[22][111] = 0;rain_draw[23][111] = 0;rain_draw[24][111] = 1;rain_draw[25][111] = 1;rain_draw[26][111] = 1;rain_draw[27][111] = 0;rain_draw[28][111] = 0;rain_draw[29][111] = 0;rain_draw[30][111] = 0;rain_draw[31][111] = 0;rain_draw[32][111] = 0;rain_draw[33][111] = 0;rain_draw[34][111] = 0;rain_draw[35][111] = 0;rain_draw[36][111] = 0;rain_draw[37][111] = 0;rain_draw[38][111] = 0;rain_draw[39][111] = 0;rain_draw[40][111] = 0;rain_draw[41][111] = 0;rain_draw[42][111] = 0;rain_draw[43][111] = 0;rain_draw[44][111] = 0;rain_draw[45][111] = 0;rain_draw[46][111] = 0;rain_draw[47][111] = 0;rain_draw[48][111] = 0;rain_draw[49][111] = 0;rain_draw[50][111] = 0;rain_draw[51][111] = 0;rain_draw[52][111] = 0;rain_draw[53][111] = 0;rain_draw[54][111] = 0;rain_draw[55][111] = 0;rain_draw[56][111] = 0;rain_draw[57][111] = 0;rain_draw[58][111] = 0;rain_draw[59][111] = 0;rain_draw[60][111] = 0;rain_draw[61][111] = 1;rain_draw[62][111] = 1;rain_draw[63][111] = 1;rain_draw[64][111] = 0;rain_draw[65][111] = 0;rain_draw[66][111] = 0;rain_draw[67][111] = 0;rain_draw[68][111] = 0;rain_draw[69][111] = 0;rain_draw[70][111] = 0;rain_draw[71][111] = 0;rain_draw[72][111] = 0;rain_draw[73][111] = 0;rain_draw[74][111] = 0;rain_draw[75][111] = 0;rain_draw[76][111] = 0;rain_draw[77][111] = 0;rain_draw[78][111] = 0;rain_draw[79][111] = 0;rain_draw[80][111] = 0;rain_draw[81][111] = 0;rain_draw[82][111] = 1;rain_draw[83][111] = 1;rain_draw[84][111] = 1;rain_draw[85][111] = 0;rain_draw[86][111] = 0;rain_draw[87][111] = 0;rain_draw[88][111] = 0;rain_draw[89][111] = 0;rain_draw[90][111] = 0;rain_draw[91][111] = 0;rain_draw[92][111] = 0;rain_draw[93][111] = 0;rain_draw[94][111] = 0;rain_draw[95][111] = 0;
        rain_draw[0][112] = 0;rain_draw[1][112] = 0;rain_draw[2][112] = 0;rain_draw[3][112] = 0;rain_draw[4][112] = 0;rain_draw[5][112] = 0;rain_draw[6][112] = 0;rain_draw[7][112] = 0;rain_draw[8][112] = 0;rain_draw[9][112] = 0;rain_draw[10][112] = 0;rain_draw[11][112] = 0;rain_draw[12][112] = 0;rain_draw[13][112] = 0;rain_draw[14][112] = 0;rain_draw[15][112] = 0;rain_draw[16][112] = 0;rain_draw[17][112] = 0;rain_draw[18][112] = 0;rain_draw[19][112] = 0;rain_draw[20][112] = 0;rain_draw[21][112] = 0;rain_draw[22][112] = 0;rain_draw[23][112] = 1;rain_draw[24][112] = 1;rain_draw[25][112] = 1;rain_draw[26][112] = 0;rain_draw[27][112] = 0;rain_draw[28][112] = 0;rain_draw[29][112] = 0;rain_draw[30][112] = 0;rain_draw[31][112] = 0;rain_draw[32][112] = 0;rain_draw[33][112] = 0;rain_draw[34][112] = 0;rain_draw[35][112] = 0;rain_draw[36][112] = 0;rain_draw[37][112] = 0;rain_draw[38][112] = 0;rain_draw[39][112] = 0;rain_draw[40][112] = 0;rain_draw[41][112] = 0;rain_draw[42][112] = 0;rain_draw[43][112] = 0;rain_draw[44][112] = 0;rain_draw[45][112] = 0;rain_draw[46][112] = 0;rain_draw[47][112] = 0;rain_draw[48][112] = 0;rain_draw[49][112] = 0;rain_draw[50][112] = 0;rain_draw[51][112] = 0;rain_draw[52][112] = 0;rain_draw[53][112] = 0;rain_draw[54][112] = 0;rain_draw[55][112] = 0;rain_draw[56][112] = 0;rain_draw[57][112] = 0;rain_draw[58][112] = 0;rain_draw[59][112] = 0;rain_draw[60][112] = 0;rain_draw[61][112] = 0;rain_draw[62][112] = 0;rain_draw[63][112] = 0;rain_draw[64][112] = 0;rain_draw[65][112] = 0;rain_draw[66][112] = 0;rain_draw[67][112] = 0;rain_draw[68][112] = 0;rain_draw[69][112] = 0;rain_draw[70][112] = 0;rain_draw[71][112] = 0;rain_draw[72][112] = 0;rain_draw[73][112] = 0;rain_draw[74][112] = 0;rain_draw[75][112] = 0;rain_draw[76][112] = 0;rain_draw[77][112] = 0;rain_draw[78][112] = 0;rain_draw[79][112] = 0;rain_draw[80][112] = 0;rain_draw[81][112] = 1;rain_draw[82][112] = 1;rain_draw[83][112] = 1;rain_draw[84][112] = 0;rain_draw[85][112] = 0;rain_draw[86][112] = 0;rain_draw[87][112] = 0;rain_draw[88][112] = 0;rain_draw[89][112] = 0;rain_draw[90][112] = 0;rain_draw[91][112] = 0;rain_draw[92][112] = 0;rain_draw[93][112] = 0;rain_draw[94][112] = 0;rain_draw[95][112] = 0;
        rain_draw[0][113] = 0;rain_draw[1][113] = 0;rain_draw[2][113] = 0;rain_draw[3][113] = 0;rain_draw[4][113] = 0;rain_draw[5][113] = 0;rain_draw[6][113] = 0;rain_draw[7][113] = 0;rain_draw[8][113] = 0;rain_draw[9][113] = 0;rain_draw[10][113] = 0;rain_draw[11][113] = 0;rain_draw[12][113] = 0;rain_draw[13][113] = 0;rain_draw[14][113] = 0;rain_draw[15][113] = 0;rain_draw[16][113] = 0;rain_draw[17][113] = 0;rain_draw[18][113] = 0;rain_draw[19][113] = 0;rain_draw[20][113] = 0;rain_draw[21][113] = 0;rain_draw[22][113] = 1;rain_draw[23][113] = 1;rain_draw[24][113] = 1;rain_draw[25][113] = 0;rain_draw[26][113] = 0;rain_draw[27][113] = 0;rain_draw[28][113] = 0;rain_draw[29][113] = 0;rain_draw[30][113] = 0;rain_draw[31][113] = 0;rain_draw[32][113] = 0;rain_draw[33][113] = 0;rain_draw[34][113] = 0;rain_draw[35][113] = 0;rain_draw[36][113] = 0;rain_draw[37][113] = 0;rain_draw[38][113] = 0;rain_draw[39][113] = 0;rain_draw[40][113] = 0;rain_draw[41][113] = 0;rain_draw[42][113] = 0;rain_draw[43][113] = 0;rain_draw[44][113] = 0;rain_draw[45][113] = 0;rain_draw[46][113] = 0;rain_draw[47][113] = 0;rain_draw[48][113] = 0;rain_draw[49][113] = 0;rain_draw[50][113] = 0;rain_draw[51][113] = 0;rain_draw[52][113] = 0;rain_draw[53][113] = 0;rain_draw[54][113] = 0;rain_draw[55][113] = 0;rain_draw[56][113] = 0;rain_draw[57][113] = 0;rain_draw[58][113] = 0;rain_draw[59][113] = 0;rain_draw[60][113] = 0;rain_draw[61][113] = 0;rain_draw[62][113] = 0;rain_draw[63][113] = 0;rain_draw[64][113] = 0;rain_draw[65][113] = 0;rain_draw[66][113] = 0;rain_draw[67][113] = 0;rain_draw[68][113] = 0;rain_draw[69][113] = 0;rain_draw[70][113] = 0;rain_draw[71][113] = 0;rain_draw[72][113] = 0;rain_draw[73][113] = 0;rain_draw[74][113] = 0;rain_draw[75][113] = 0;rain_draw[76][113] = 0;rain_draw[77][113] = 0;rain_draw[78][113] = 0;rain_draw[79][113] = 0;rain_draw[80][113] = 1;rain_draw[81][113] = 1;rain_draw[82][113] = 1;rain_draw[83][113] = 0;rain_draw[84][113] = 0;rain_draw[85][113] = 0;rain_draw[86][113] = 0;rain_draw[87][113] = 0;rain_draw[88][113] = 0;rain_draw[89][113] = 0;rain_draw[90][113] = 0;rain_draw[91][113] = 0;rain_draw[92][113] = 0;rain_draw[93][113] = 0;rain_draw[94][113] = 0;rain_draw[95][113] = 0;
        rain_draw[0][114] = 0;rain_draw[1][114] = 0;rain_draw[2][114] = 0;rain_draw[3][114] = 0;rain_draw[4][114] = 0;rain_draw[5][114] = 0;rain_draw[6][114] = 0;rain_draw[7][114] = 0;rain_draw[8][114] = 0;rain_draw[9][114] = 0;rain_draw[10][114] = 0;rain_draw[11][114] = 0;rain_draw[12][114] = 0;rain_draw[13][114] = 0;rain_draw[14][114] = 0;rain_draw[15][114] = 0;rain_draw[16][114] = 0;rain_draw[17][114] = 0;rain_draw[18][114] = 0;rain_draw[19][114] = 0;rain_draw[20][114] = 0;rain_draw[21][114] = 1;rain_draw[22][114] = 1;rain_draw[23][114] = 1;rain_draw[24][114] = 0;rain_draw[25][114] = 0;rain_draw[26][114] = 0;rain_draw[27][114] = 0;rain_draw[28][114] = 0;rain_draw[29][114] = 0;rain_draw[30][114] = 0;rain_draw[31][114] = 0;rain_draw[32][114] = 0;rain_draw[33][114] = 0;rain_draw[34][114] = 0;rain_draw[35][114] = 0;rain_draw[36][114] = 0;rain_draw[37][114] = 0;rain_draw[38][114] = 0;rain_draw[39][114] = 0;rain_draw[40][114] = 0;rain_draw[41][114] = 0;rain_draw[42][114] = 0;rain_draw[43][114] = 0;rain_draw[44][114] = 0;rain_draw[45][114] = 0;rain_draw[46][114] = 0;rain_draw[47][114] = 0;rain_draw[48][114] = 0;rain_draw[49][114] = 0;rain_draw[50][114] = 0;rain_draw[51][114] = 0;rain_draw[52][114] = 0;rain_draw[53][114] = 0;rain_draw[54][114] = 0;rain_draw[55][114] = 0;rain_draw[56][114] = 0;rain_draw[57][114] = 0;rain_draw[58][114] = 0;rain_draw[59][114] = 0;rain_draw[60][114] = 0;rain_draw[61][114] = 0;rain_draw[62][114] = 0;rain_draw[63][114] = 0;rain_draw[64][114] = 0;rain_draw[65][114] = 0;rain_draw[66][114] = 0;rain_draw[67][114] = 0;rain_draw[68][114] = 0;rain_draw[69][114] = 0;rain_draw[70][114] = 0;rain_draw[71][114] = 0;rain_draw[72][114] = 0;rain_draw[73][114] = 0;rain_draw[74][114] = 0;rain_draw[75][114] = 0;rain_draw[76][114] = 0;rain_draw[77][114] = 0;rain_draw[78][114] = 0;rain_draw[79][114] = 0;rain_draw[80][114] = 0;rain_draw[81][114] = 0;rain_draw[82][114] = 0;rain_draw[83][114] = 0;rain_draw[84][114] = 0;rain_draw[85][114] = 0;rain_draw[86][114] = 0;rain_draw[87][114] = 0;rain_draw[88][114] = 0;rain_draw[89][114] = 0;rain_draw[90][114] = 0;rain_draw[91][114] = 0;rain_draw[92][114] = 0;rain_draw[93][114] = 0;rain_draw[94][114] = 0;rain_draw[95][114] = 0;
        rain_draw[0][115] = 0;rain_draw[1][115] = 0;rain_draw[2][115] = 0;rain_draw[3][115] = 0;rain_draw[4][115] = 0;rain_draw[5][115] = 0;rain_draw[6][115] = 0;rain_draw[7][115] = 0;rain_draw[8][115] = 0;rain_draw[9][115] = 0;rain_draw[10][115] = 0;rain_draw[11][115] = 0;rain_draw[12][115] = 0;rain_draw[13][115] = 0;rain_draw[14][115] = 0;rain_draw[15][115] = 0;rain_draw[16][115] = 0;rain_draw[17][115] = 0;rain_draw[18][115] = 0;rain_draw[19][115] = 0;rain_draw[20][115] = 0;rain_draw[21][115] = 0;rain_draw[22][115] = 0;rain_draw[23][115] = 0;rain_draw[24][115] = 0;rain_draw[25][115] = 0;rain_draw[26][115] = 0;rain_draw[27][115] = 0;rain_draw[28][115] = 0;rain_draw[29][115] = 0;rain_draw[30][115] = 0;rain_draw[31][115] = 0;rain_draw[32][115] = 0;rain_draw[33][115] = 0;rain_draw[34][115] = 0;rain_draw[35][115] = 0;rain_draw[36][115] = 0;rain_draw[37][115] = 0;rain_draw[38][115] = 0;rain_draw[39][115] = 0;rain_draw[40][115] = 0;rain_draw[41][115] = 0;rain_draw[42][115] = 0;rain_draw[43][115] = 0;rain_draw[44][115] = 0;rain_draw[45][115] = 0;rain_draw[46][115] = 0;rain_draw[47][115] = 0;rain_draw[48][115] = 0;rain_draw[49][115] = 0;rain_draw[50][115] = 0;rain_draw[51][115] = 0;rain_draw[52][115] = 0;rain_draw[53][115] = 0;rain_draw[54][115] = 0;rain_draw[55][115] = 0;rain_draw[56][115] = 0;rain_draw[57][115] = 0;rain_draw[58][115] = 0;rain_draw[59][115] = 0;rain_draw[60][115] = 0;rain_draw[61][115] = 0;rain_draw[62][115] = 0;rain_draw[63][115] = 0;rain_draw[64][115] = 0;rain_draw[65][115] = 0;rain_draw[66][115] = 0;rain_draw[67][115] = 0;rain_draw[68][115] = 0;rain_draw[69][115] = 0;rain_draw[70][115] = 0;rain_draw[71][115] = 0;rain_draw[72][115] = 0;rain_draw[73][115] = 0;rain_draw[74][115] = 0;rain_draw[75][115] = 0;rain_draw[76][115] = 0;rain_draw[77][115] = 0;rain_draw[78][115] = 0;rain_draw[79][115] = 0;rain_draw[80][115] = 0;rain_draw[81][115] = 0;rain_draw[82][115] = 0;rain_draw[83][115] = 0;rain_draw[84][115] = 0;rain_draw[85][115] = 0;rain_draw[86][115] = 0;rain_draw[87][115] = 0;rain_draw[88][115] = 0;rain_draw[89][115] = 0;rain_draw[90][115] = 0;rain_draw[91][115] = 0;rain_draw[92][115] = 0;rain_draw[93][115] = 0;rain_draw[94][115] = 0;rain_draw[95][115] = 0;
        rain_draw[0][116] = 0;rain_draw[1][116] = 0;rain_draw[2][116] = 0;rain_draw[3][116] = 0;rain_draw[4][116] = 0;rain_draw[5][116] = 0;rain_draw[6][116] = 0;rain_draw[7][116] = 0;rain_draw[8][116] = 0;rain_draw[9][116] = 0;rain_draw[10][116] = 0;rain_draw[11][116] = 0;rain_draw[12][116] = 0;rain_draw[13][116] = 0;rain_draw[14][116] = 0;rain_draw[15][116] = 0;rain_draw[16][116] = 0;rain_draw[17][116] = 0;rain_draw[18][116] = 0;rain_draw[19][116] = 0;rain_draw[20][116] = 0;rain_draw[21][116] = 0;rain_draw[22][116] = 0;rain_draw[23][116] = 0;rain_draw[24][116] = 0;rain_draw[25][116] = 0;rain_draw[26][116] = 0;rain_draw[27][116] = 0;rain_draw[28][116] = 0;rain_draw[29][116] = 0;rain_draw[30][116] = 0;rain_draw[31][116] = 0;rain_draw[32][116] = 0;rain_draw[33][116] = 0;rain_draw[34][116] = 0;rain_draw[35][116] = 0;rain_draw[36][116] = 0;rain_draw[37][116] = 0;rain_draw[38][116] = 0;rain_draw[39][116] = 0;rain_draw[40][116] = 0;rain_draw[41][116] = 0;rain_draw[42][116] = 0;rain_draw[43][116] = 0;rain_draw[44][116] = 0;rain_draw[45][116] = 0;rain_draw[46][116] = 0;rain_draw[47][116] = 0;rain_draw[48][116] = 0;rain_draw[49][116] = 0;rain_draw[50][116] = 0;rain_draw[51][116] = 0;rain_draw[52][116] = 0;rain_draw[53][116] = 0;rain_draw[54][116] = 0;rain_draw[55][116] = 0;rain_draw[56][116] = 0;rain_draw[57][116] = 0;rain_draw[58][116] = 0;rain_draw[59][116] = 0;rain_draw[60][116] = 0;rain_draw[61][116] = 0;rain_draw[62][116] = 0;rain_draw[63][116] = 0;rain_draw[64][116] = 0;rain_draw[65][116] = 0;rain_draw[66][116] = 0;rain_draw[67][116] = 0;rain_draw[68][116] = 0;rain_draw[69][116] = 0;rain_draw[70][116] = 0;rain_draw[71][116] = 0;rain_draw[72][116] = 0;rain_draw[73][116] = 0;rain_draw[74][116] = 0;rain_draw[75][116] = 0;rain_draw[76][116] = 0;rain_draw[77][116] = 0;rain_draw[78][116] = 0;rain_draw[79][116] = 0;rain_draw[80][116] = 0;rain_draw[81][116] = 0;rain_draw[82][116] = 0;rain_draw[83][116] = 0;rain_draw[84][116] = 0;rain_draw[85][116] = 0;rain_draw[86][116] = 0;rain_draw[87][116] = 0;rain_draw[88][116] = 0;rain_draw[89][116] = 0;rain_draw[90][116] = 0;rain_draw[91][116] = 0;rain_draw[92][116] = 0;rain_draw[93][116] = 0;rain_draw[94][116] = 0;rain_draw[95][116] = 0;
        rain_draw[0][117] = 0;rain_draw[1][117] = 0;rain_draw[2][117] = 0;rain_draw[3][117] = 0;rain_draw[4][117] = 0;rain_draw[5][117] = 0;rain_draw[6][117] = 0;rain_draw[7][117] = 0;rain_draw[8][117] = 0;rain_draw[9][117] = 0;rain_draw[10][117] = 0;rain_draw[11][117] = 0;rain_draw[12][117] = 0;rain_draw[13][117] = 0;rain_draw[14][117] = 0;rain_draw[15][117] = 0;rain_draw[16][117] = 0;rain_draw[17][117] = 0;rain_draw[18][117] = 0;rain_draw[19][117] = 0;rain_draw[20][117] = 0;rain_draw[21][117] = 0;rain_draw[22][117] = 0;rain_draw[23][117] = 0;rain_draw[24][117] = 0;rain_draw[25][117] = 0;rain_draw[26][117] = 0;rain_draw[27][117] = 0;rain_draw[28][117] = 0;rain_draw[29][117] = 0;rain_draw[30][117] = 0;rain_draw[31][117] = 0;rain_draw[32][117] = 0;rain_draw[33][117] = 0;rain_draw[34][117] = 0;rain_draw[35][117] = 0;rain_draw[36][117] = 0;rain_draw[37][117] = 0;rain_draw[38][117] = 0;rain_draw[39][117] = 0;rain_draw[40][117] = 0;rain_draw[41][117] = 0;rain_draw[42][117] = 0;rain_draw[43][117] = 0;rain_draw[44][117] = 0;rain_draw[45][117] = 0;rain_draw[46][117] = 0;rain_draw[47][117] = 0;rain_draw[48][117] = 0;rain_draw[49][117] = 0;rain_draw[50][117] = 1;rain_draw[51][117] = 1;rain_draw[52][117] = 1;rain_draw[53][117] = 0;rain_draw[54][117] = 0;rain_draw[55][117] = 0;rain_draw[56][117] = 0;rain_draw[57][117] = 0;rain_draw[58][117] = 0;rain_draw[59][117] = 0;rain_draw[60][117] = 0;rain_draw[61][117] = 0;rain_draw[62][117] = 0;rain_draw[63][117] = 0;rain_draw[64][117] = 0;rain_draw[65][117] = 0;rain_draw[66][117] = 0;rain_draw[67][117] = 0;rain_draw[68][117] = 0;rain_draw[69][117] = 0;rain_draw[70][117] = 0;rain_draw[71][117] = 0;rain_draw[72][117] = 0;rain_draw[73][117] = 0;rain_draw[74][117] = 0;rain_draw[75][117] = 0;rain_draw[76][117] = 0;rain_draw[77][117] = 0;rain_draw[78][117] = 0;rain_draw[79][117] = 0;rain_draw[80][117] = 0;rain_draw[81][117] = 0;rain_draw[82][117] = 0;rain_draw[83][117] = 0;rain_draw[84][117] = 0;rain_draw[85][117] = 0;rain_draw[86][117] = 0;rain_draw[87][117] = 0;rain_draw[88][117] = 0;rain_draw[89][117] = 0;rain_draw[90][117] = 0;rain_draw[91][117] = 0;rain_draw[92][117] = 0;rain_draw[93][117] = 0;rain_draw[94][117] = 0;rain_draw[95][117] = 0;
        rain_draw[0][118] = 0;rain_draw[1][118] = 0;rain_draw[2][118] = 0;rain_draw[3][118] = 0;rain_draw[4][118] = 0;rain_draw[5][118] = 0;rain_draw[6][118] = 0;rain_draw[7][118] = 0;rain_draw[8][118] = 0;rain_draw[9][118] = 0;rain_draw[10][118] = 0;rain_draw[11][118] = 0;rain_draw[12][118] = 0;rain_draw[13][118] = 0;rain_draw[14][118] = 0;rain_draw[15][118] = 0;rain_draw[16][118] = 0;rain_draw[17][118] = 0;rain_draw[18][118] = 0;rain_draw[19][118] = 0;rain_draw[20][118] = 0;rain_draw[21][118] = 0;rain_draw[22][118] = 0;rain_draw[23][118] = 0;rain_draw[24][118] = 0;rain_draw[25][118] = 0;rain_draw[26][118] = 0;rain_draw[27][118] = 0;rain_draw[28][118] = 0;rain_draw[29][118] = 0;rain_draw[30][118] = 0;rain_draw[31][118] = 0;rain_draw[32][118] = 0;rain_draw[33][118] = 0;rain_draw[34][118] = 0;rain_draw[35][118] = 0;rain_draw[36][118] = 0;rain_draw[37][118] = 0;rain_draw[38][118] = 0;rain_draw[39][118] = 0;rain_draw[40][118] = 0;rain_draw[41][118] = 0;rain_draw[42][118] = 0;rain_draw[43][118] = 0;rain_draw[44][118] = 0;rain_draw[45][118] = 0;rain_draw[46][118] = 0;rain_draw[47][118] = 0;rain_draw[48][118] = 0;rain_draw[49][118] = 1;rain_draw[50][118] = 1;rain_draw[51][118] = 1;rain_draw[52][118] = 0;rain_draw[53][118] = 0;rain_draw[54][118] = 0;rain_draw[55][118] = 0;rain_draw[56][118] = 0;rain_draw[57][118] = 0;rain_draw[58][118] = 0;rain_draw[59][118] = 0;rain_draw[60][118] = 0;rain_draw[61][118] = 0;rain_draw[62][118] = 0;rain_draw[63][118] = 0;rain_draw[64][118] = 0;rain_draw[65][118] = 0;rain_draw[66][118] = 0;rain_draw[67][118] = 0;rain_draw[68][118] = 0;rain_draw[69][118] = 0;rain_draw[70][118] = 0;rain_draw[71][118] = 0;rain_draw[72][118] = 0;rain_draw[73][118] = 0;rain_draw[74][118] = 0;rain_draw[75][118] = 0;rain_draw[76][118] = 0;rain_draw[77][118] = 0;rain_draw[78][118] = 0;rain_draw[79][118] = 0;rain_draw[80][118] = 0;rain_draw[81][118] = 0;rain_draw[82][118] = 0;rain_draw[83][118] = 0;rain_draw[84][118] = 0;rain_draw[85][118] = 0;rain_draw[86][118] = 0;rain_draw[87][118] = 0;rain_draw[88][118] = 0;rain_draw[89][118] = 0;rain_draw[90][118] = 0;rain_draw[91][118] = 0;rain_draw[92][118] = 0;rain_draw[93][118] = 0;rain_draw[94][118] = 0;rain_draw[95][118] = 0;
        rain_draw[0][119] = 0;rain_draw[1][119] = 0;rain_draw[2][119] = 0;rain_draw[3][119] = 0;rain_draw[4][119] = 0;rain_draw[5][119] = 0;rain_draw[6][119] = 0;rain_draw[7][119] = 0;rain_draw[8][119] = 0;rain_draw[9][119] = 0;rain_draw[10][119] = 0;rain_draw[11][119] = 0;rain_draw[12][119] = 0;rain_draw[13][119] = 0;rain_draw[14][119] = 0;rain_draw[15][119] = 0;rain_draw[16][119] = 0;rain_draw[17][119] = 0;rain_draw[18][119] = 0;rain_draw[19][119] = 0;rain_draw[20][119] = 0;rain_draw[21][119] = 0;rain_draw[22][119] = 0;rain_draw[23][119] = 0;rain_draw[24][119] = 0;rain_draw[25][119] = 0;rain_draw[26][119] = 0;rain_draw[27][119] = 0;rain_draw[28][119] = 0;rain_draw[29][119] = 0;rain_draw[30][119] = 0;rain_draw[31][119] = 0;rain_draw[32][119] = 0;rain_draw[33][119] = 0;rain_draw[34][119] = 0;rain_draw[35][119] = 0;rain_draw[36][119] = 0;rain_draw[37][119] = 0;rain_draw[38][119] = 0;rain_draw[39][119] = 0;rain_draw[40][119] = 0;rain_draw[41][119] = 0;rain_draw[42][119] = 0;rain_draw[43][119] = 0;rain_draw[44][119] = 0;rain_draw[45][119] = 0;rain_draw[46][119] = 0;rain_draw[47][119] = 0;rain_draw[48][119] = 1;rain_draw[49][119] = 1;rain_draw[50][119] = 1;rain_draw[51][119] = 0;rain_draw[52][119] = 0;rain_draw[53][119] = 0;rain_draw[54][119] = 0;rain_draw[55][119] = 0;rain_draw[56][119] = 0;rain_draw[57][119] = 0;rain_draw[58][119] = 0;rain_draw[59][119] = 0;rain_draw[60][119] = 0;rain_draw[61][119] = 0;rain_draw[62][119] = 0;rain_draw[63][119] = 0;rain_draw[64][119] = 0;rain_draw[65][119] = 0;rain_draw[66][119] = 0;rain_draw[67][119] = 0;rain_draw[68][119] = 0;rain_draw[69][119] = 0;rain_draw[70][119] = 0;rain_draw[71][119] = 0;rain_draw[72][119] = 0;rain_draw[73][119] = 0;rain_draw[74][119] = 0;rain_draw[75][119] = 0;rain_draw[76][119] = 0;rain_draw[77][119] = 0;rain_draw[78][119] = 0;rain_draw[79][119] = 0;rain_draw[80][119] = 0;rain_draw[81][119] = 0;rain_draw[82][119] = 0;rain_draw[83][119] = 0;rain_draw[84][119] = 0;rain_draw[85][119] = 0;rain_draw[86][119] = 0;rain_draw[87][119] = 0;rain_draw[88][119] = 0;rain_draw[89][119] = 0;rain_draw[90][119] = 0;rain_draw[91][119] = 0;rain_draw[92][119] = 0;rain_draw[93][119] = 0;rain_draw[94][119] = 0;rain_draw[95][119] = 0;
        rain_draw[0][120] = 0;rain_draw[1][120] = 0;rain_draw[2][120] = 0;rain_draw[3][120] = 0;rain_draw[4][120] = 0;rain_draw[5][120] = 0;rain_draw[6][120] = 0;rain_draw[7][120] = 0;rain_draw[8][120] = 0;rain_draw[9][120] = 0;rain_draw[10][120] = 0;rain_draw[11][120] = 0;rain_draw[12][120] = 0;rain_draw[13][120] = 0;rain_draw[14][120] = 0;rain_draw[15][120] = 0;rain_draw[16][120] = 0;rain_draw[17][120] = 0;rain_draw[18][120] = 0;rain_draw[19][120] = 0;rain_draw[20][120] = 0;rain_draw[21][120] = 0;rain_draw[22][120] = 0;rain_draw[23][120] = 0;rain_draw[24][120] = 0;rain_draw[25][120] = 0;rain_draw[26][120] = 0;rain_draw[27][120] = 0;rain_draw[28][120] = 0;rain_draw[29][120] = 0;rain_draw[30][120] = 0;rain_draw[31][120] = 0;rain_draw[32][120] = 0;rain_draw[33][120] = 0;rain_draw[34][120] = 0;rain_draw[35][120] = 0;rain_draw[36][120] = 0;rain_draw[37][120] = 0;rain_draw[38][120] = 0;rain_draw[39][120] = 0;rain_draw[40][120] = 0;rain_draw[41][120] = 0;rain_draw[42][120] = 0;rain_draw[43][120] = 0;rain_draw[44][120] = 0;rain_draw[45][120] = 0;rain_draw[46][120] = 0;rain_draw[47][120] = 1;rain_draw[48][120] = 1;rain_draw[49][120] = 1;rain_draw[50][120] = 0;rain_draw[51][120] = 0;rain_draw[52][120] = 0;rain_draw[53][120] = 0;rain_draw[54][120] = 0;rain_draw[55][120] = 0;rain_draw[56][120] = 0;rain_draw[57][120] = 0;rain_draw[58][120] = 0;rain_draw[59][120] = 0;rain_draw[60][120] = 0;rain_draw[61][120] = 0;rain_draw[62][120] = 0;rain_draw[63][120] = 0;rain_draw[64][120] = 0;rain_draw[65][120] = 0;rain_draw[66][120] = 0;rain_draw[67][120] = 0;rain_draw[68][120] = 0;rain_draw[69][120] = 0;rain_draw[70][120] = 0;rain_draw[71][120] = 0;rain_draw[72][120] = 0;rain_draw[73][120] = 0;rain_draw[74][120] = 0;rain_draw[75][120] = 0;rain_draw[76][120] = 0;rain_draw[77][120] = 0;rain_draw[78][120] = 0;rain_draw[79][120] = 0;rain_draw[80][120] = 0;rain_draw[81][120] = 0;rain_draw[82][120] = 0;rain_draw[83][120] = 0;rain_draw[84][120] = 0;rain_draw[85][120] = 0;rain_draw[86][120] = 0;rain_draw[87][120] = 0;rain_draw[88][120] = 0;rain_draw[89][120] = 0;rain_draw[90][120] = 0;rain_draw[91][120] = 0;rain_draw[92][120] = 0;rain_draw[93][120] = 0;rain_draw[94][120] = 0;rain_draw[95][120] = 0;
        rain_draw[0][121] = 0;rain_draw[1][121] = 0;rain_draw[2][121] = 0;rain_draw[3][121] = 0;rain_draw[4][121] = 0;rain_draw[5][121] = 0;rain_draw[6][121] = 0;rain_draw[7][121] = 0;rain_draw[8][121] = 0;rain_draw[9][121] = 0;rain_draw[10][121] = 0;rain_draw[11][121] = 0;rain_draw[12][121] = 0;rain_draw[13][121] = 0;rain_draw[14][121] = 0;rain_draw[15][121] = 0;rain_draw[16][121] = 0;rain_draw[17][121] = 0;rain_draw[18][121] = 0;rain_draw[19][121] = 0;rain_draw[20][121] = 0;rain_draw[21][121] = 0;rain_draw[22][121] = 0;rain_draw[23][121] = 0;rain_draw[24][121] = 0;rain_draw[25][121] = 0;rain_draw[26][121] = 0;rain_draw[27][121] = 0;rain_draw[28][121] = 0;rain_draw[29][121] = 0;rain_draw[30][121] = 0;rain_draw[31][121] = 0;rain_draw[32][121] = 0;rain_draw[33][121] = 0;rain_draw[34][121] = 0;rain_draw[35][121] = 0;rain_draw[36][121] = 0;rain_draw[37][121] = 0;rain_draw[38][121] = 0;rain_draw[39][121] = 0;rain_draw[40][121] = 0;rain_draw[41][121] = 0;rain_draw[42][121] = 0;rain_draw[43][121] = 0;rain_draw[44][121] = 0;rain_draw[45][121] = 0;rain_draw[46][121] = 1;rain_draw[47][121] = 1;rain_draw[48][121] = 1;rain_draw[49][121] = 0;rain_draw[50][121] = 0;rain_draw[51][121] = 0;rain_draw[52][121] = 0;rain_draw[53][121] = 0;rain_draw[54][121] = 0;rain_draw[55][121] = 0;rain_draw[56][121] = 0;rain_draw[57][121] = 0;rain_draw[58][121] = 0;rain_draw[59][121] = 0;rain_draw[60][121] = 0;rain_draw[61][121] = 0;rain_draw[62][121] = 0;rain_draw[63][121] = 0;rain_draw[64][121] = 0;rain_draw[65][121] = 0;rain_draw[66][121] = 0;rain_draw[67][121] = 0;rain_draw[68][121] = 0;rain_draw[69][121] = 0;rain_draw[70][121] = 0;rain_draw[71][121] = 0;rain_draw[72][121] = 0;rain_draw[73][121] = 0;rain_draw[74][121] = 0;rain_draw[75][121] = 0;rain_draw[76][121] = 0;rain_draw[77][121] = 0;rain_draw[78][121] = 0;rain_draw[79][121] = 0;rain_draw[80][121] = 0;rain_draw[81][121] = 0;rain_draw[82][121] = 0;rain_draw[83][121] = 0;rain_draw[84][121] = 0;rain_draw[85][121] = 0;rain_draw[86][121] = 0;rain_draw[87][121] = 0;rain_draw[88][121] = 0;rain_draw[89][121] = 0;rain_draw[90][121] = 0;rain_draw[91][121] = 0;rain_draw[92][121] = 0;rain_draw[93][121] = 0;rain_draw[94][121] = 0;rain_draw[95][121] = 0;
        rain_draw[0][122] = 0;rain_draw[1][122] = 0;rain_draw[2][122] = 0;rain_draw[3][122] = 0;rain_draw[4][122] = 0;rain_draw[5][122] = 0;rain_draw[6][122] = 0;rain_draw[7][122] = 0;rain_draw[8][122] = 0;rain_draw[9][122] = 0;rain_draw[10][122] = 0;rain_draw[11][122] = 0;rain_draw[12][122] = 0;rain_draw[13][122] = 0;rain_draw[14][122] = 0;rain_draw[15][122] = 0;rain_draw[16][122] = 0;rain_draw[17][122] = 0;rain_draw[18][122] = 0;rain_draw[19][122] = 0;rain_draw[20][122] = 0;rain_draw[21][122] = 0;rain_draw[22][122] = 0;rain_draw[23][122] = 0;rain_draw[24][122] = 0;rain_draw[25][122] = 0;rain_draw[26][122] = 0;rain_draw[27][122] = 0;rain_draw[28][122] = 0;rain_draw[29][122] = 0;rain_draw[30][122] = 0;rain_draw[31][122] = 0;rain_draw[32][122] = 0;rain_draw[33][122] = 0;rain_draw[34][122] = 0;rain_draw[35][122] = 0;rain_draw[36][122] = 0;rain_draw[37][122] = 0;rain_draw[38][122] = 0;rain_draw[39][122] = 0;rain_draw[40][122] = 0;rain_draw[41][122] = 0;rain_draw[42][122] = 0;rain_draw[43][122] = 0;rain_draw[44][122] = 0;rain_draw[45][122] = 1;rain_draw[46][122] = 1;rain_draw[47][122] = 1;rain_draw[48][122] = 0;rain_draw[49][122] = 0;rain_draw[50][122] = 0;rain_draw[51][122] = 0;rain_draw[52][122] = 0;rain_draw[53][122] = 0;rain_draw[54][122] = 0;rain_draw[55][122] = 0;rain_draw[56][122] = 0;rain_draw[57][122] = 0;rain_draw[58][122] = 0;rain_draw[59][122] = 0;rain_draw[60][122] = 0;rain_draw[61][122] = 0;rain_draw[62][122] = 0;rain_draw[63][122] = 0;rain_draw[64][122] = 0;rain_draw[65][122] = 0;rain_draw[66][122] = 0;rain_draw[67][122] = 0;rain_draw[68][122] = 0;rain_draw[69][122] = 0;rain_draw[70][122] = 0;rain_draw[71][122] = 0;rain_draw[72][122] = 0;rain_draw[73][122] = 0;rain_draw[74][122] = 0;rain_draw[75][122] = 0;rain_draw[76][122] = 0;rain_draw[77][122] = 0;rain_draw[78][122] = 0;rain_draw[79][122] = 0;rain_draw[80][122] = 0;rain_draw[81][122] = 0;rain_draw[82][122] = 0;rain_draw[83][122] = 0;rain_draw[84][122] = 0;rain_draw[85][122] = 0;rain_draw[86][122] = 0;rain_draw[87][122] = 0;rain_draw[88][122] = 0;rain_draw[89][122] = 0;rain_draw[90][122] = 0;rain_draw[91][122] = 0;rain_draw[92][122] = 0;rain_draw[93][122] = 0;rain_draw[94][122] = 0;rain_draw[95][122] = 0;
        rain_draw[0][123] = 0;rain_draw[1][123] = 0;rain_draw[2][123] = 0;rain_draw[3][123] = 0;rain_draw[4][123] = 0;rain_draw[5][123] = 0;rain_draw[6][123] = 0;rain_draw[7][123] = 0;rain_draw[8][123] = 0;rain_draw[9][123] = 0;rain_draw[10][123] = 0;rain_draw[11][123] = 0;rain_draw[12][123] = 0;rain_draw[13][123] = 0;rain_draw[14][123] = 0;rain_draw[15][123] = 0;rain_draw[16][123] = 0;rain_draw[17][123] = 0;rain_draw[18][123] = 0;rain_draw[19][123] = 0;rain_draw[20][123] = 0;rain_draw[21][123] = 0;rain_draw[22][123] = 0;rain_draw[23][123] = 0;rain_draw[24][123] = 0;rain_draw[25][123] = 0;rain_draw[26][123] = 0;rain_draw[27][123] = 0;rain_draw[28][123] = 0;rain_draw[29][123] = 0;rain_draw[30][123] = 0;rain_draw[31][123] = 0;rain_draw[32][123] = 0;rain_draw[33][123] = 0;rain_draw[34][123] = 0;rain_draw[35][123] = 0;rain_draw[36][123] = 0;rain_draw[37][123] = 0;rain_draw[38][123] = 0;rain_draw[39][123] = 0;rain_draw[40][123] = 0;rain_draw[41][123] = 0;rain_draw[42][123] = 0;rain_draw[43][123] = 0;rain_draw[44][123] = 1;rain_draw[45][123] = 1;rain_draw[46][123] = 1;rain_draw[47][123] = 0;rain_draw[48][123] = 0;rain_draw[49][123] = 0;rain_draw[50][123] = 0;rain_draw[51][123] = 0;rain_draw[52][123] = 0;rain_draw[53][123] = 0;rain_draw[54][123] = 0;rain_draw[55][123] = 0;rain_draw[56][123] = 0;rain_draw[57][123] = 0;rain_draw[58][123] = 0;rain_draw[59][123] = 0;rain_draw[60][123] = 0;rain_draw[61][123] = 0;rain_draw[62][123] = 0;rain_draw[63][123] = 0;rain_draw[64][123] = 0;rain_draw[65][123] = 0;rain_draw[66][123] = 0;rain_draw[67][123] = 0;rain_draw[68][123] = 0;rain_draw[69][123] = 0;rain_draw[70][123] = 0;rain_draw[71][123] = 0;rain_draw[72][123] = 0;rain_draw[73][123] = 0;rain_draw[74][123] = 0;rain_draw[75][123] = 0;rain_draw[76][123] = 0;rain_draw[77][123] = 0;rain_draw[78][123] = 0;rain_draw[79][123] = 0;rain_draw[80][123] = 0;rain_draw[81][123] = 0;rain_draw[82][123] = 0;rain_draw[83][123] = 0;rain_draw[84][123] = 0;rain_draw[85][123] = 0;rain_draw[86][123] = 0;rain_draw[87][123] = 0;rain_draw[88][123] = 0;rain_draw[89][123] = 0;rain_draw[90][123] = 0;rain_draw[91][123] = 0;rain_draw[92][123] = 0;rain_draw[93][123] = 0;rain_draw[94][123] = 0;rain_draw[95][123] = 0;
        rain_draw[0][124] = 0;rain_draw[1][124] = 0;rain_draw[2][124] = 0;rain_draw[3][124] = 0;rain_draw[4][124] = 0;rain_draw[5][124] = 0;rain_draw[6][124] = 0;rain_draw[7][124] = 0;rain_draw[8][124] = 0;rain_draw[9][124] = 0;rain_draw[10][124] = 0;rain_draw[11][124] = 0;rain_draw[12][124] = 0;rain_draw[13][124] = 0;rain_draw[14][124] = 0;rain_draw[15][124] = 0;rain_draw[16][124] = 0;rain_draw[17][124] = 0;rain_draw[18][124] = 0;rain_draw[19][124] = 0;rain_draw[20][124] = 0;rain_draw[21][124] = 0;rain_draw[22][124] = 0;rain_draw[23][124] = 0;rain_draw[24][124] = 0;rain_draw[25][124] = 0;rain_draw[26][124] = 0;rain_draw[27][124] = 0;rain_draw[28][124] = 0;rain_draw[29][124] = 0;rain_draw[30][124] = 0;rain_draw[31][124] = 0;rain_draw[32][124] = 0;rain_draw[33][124] = 0;rain_draw[34][124] = 0;rain_draw[35][124] = 0;rain_draw[36][124] = 0;rain_draw[37][124] = 0;rain_draw[38][124] = 0;rain_draw[39][124] = 0;rain_draw[40][124] = 0;rain_draw[41][124] = 0;rain_draw[42][124] = 0;rain_draw[43][124] = 0;rain_draw[44][124] = 0;rain_draw[45][124] = 0;rain_draw[46][124] = 0;rain_draw[47][124] = 0;rain_draw[48][124] = 0;rain_draw[49][124] = 0;rain_draw[50][124] = 0;rain_draw[51][124] = 0;rain_draw[52][124] = 0;rain_draw[53][124] = 0;rain_draw[54][124] = 0;rain_draw[55][124] = 0;rain_draw[56][124] = 0;rain_draw[57][124] = 0;rain_draw[58][124] = 0;rain_draw[59][124] = 0;rain_draw[60][124] = 0;rain_draw[61][124] = 0;rain_draw[62][124] = 0;rain_draw[63][124] = 0;rain_draw[64][124] = 0;rain_draw[65][124] = 0;rain_draw[66][124] = 0;rain_draw[67][124] = 0;rain_draw[68][124] = 0;rain_draw[69][124] = 0;rain_draw[70][124] = 0;rain_draw[71][124] = 0;rain_draw[72][124] = 0;rain_draw[73][124] = 0;rain_draw[74][124] = 0;rain_draw[75][124] = 0;rain_draw[76][124] = 0;rain_draw[77][124] = 0;rain_draw[78][124] = 0;rain_draw[79][124] = 0;rain_draw[80][124] = 0;rain_draw[81][124] = 0;rain_draw[82][124] = 0;rain_draw[83][124] = 0;rain_draw[84][124] = 0;rain_draw[85][124] = 0;rain_draw[86][124] = 0;rain_draw[87][124] = 0;rain_draw[88][124] = 0;rain_draw[89][124] = 0;rain_draw[90][124] = 0;rain_draw[91][124] = 0;rain_draw[92][124] = 0;rain_draw[93][124] = 0;rain_draw[94][124] = 0;rain_draw[95][124] = 0;
        rain_draw[0][125] = 0;rain_draw[1][125] = 0;rain_draw[2][125] = 0;rain_draw[3][125] = 0;rain_draw[4][125] = 0;rain_draw[5][125] = 0;rain_draw[6][125] = 0;rain_draw[7][125] = 0;rain_draw[8][125] = 0;rain_draw[9][125] = 0;rain_draw[10][125] = 0;rain_draw[11][125] = 0;rain_draw[12][125] = 0;rain_draw[13][125] = 0;rain_draw[14][125] = 0;rain_draw[15][125] = 0;rain_draw[16][125] = 0;rain_draw[17][125] = 0;rain_draw[18][125] = 0;rain_draw[19][125] = 0;rain_draw[20][125] = 0;rain_draw[21][125] = 0;rain_draw[22][125] = 0;rain_draw[23][125] = 0;rain_draw[24][125] = 0;rain_draw[25][125] = 0;rain_draw[26][125] = 0;rain_draw[27][125] = 0;rain_draw[28][125] = 0;rain_draw[29][125] = 0;rain_draw[30][125] = 0;rain_draw[31][125] = 0;rain_draw[32][125] = 0;rain_draw[33][125] = 0;rain_draw[34][125] = 0;rain_draw[35][125] = 0;rain_draw[36][125] = 0;rain_draw[37][125] = 0;rain_draw[38][125] = 0;rain_draw[39][125] = 0;rain_draw[40][125] = 0;rain_draw[41][125] = 0;rain_draw[42][125] = 0;rain_draw[43][125] = 0;rain_draw[44][125] = 0;rain_draw[45][125] = 0;rain_draw[46][125] = 0;rain_draw[47][125] = 0;rain_draw[48][125] = 0;rain_draw[49][125] = 0;rain_draw[50][125] = 0;rain_draw[51][125] = 0;rain_draw[52][125] = 0;rain_draw[53][125] = 0;rain_draw[54][125] = 0;rain_draw[55][125] = 0;rain_draw[56][125] = 0;rain_draw[57][125] = 0;rain_draw[58][125] = 0;rain_draw[59][125] = 0;rain_draw[60][125] = 0;rain_draw[61][125] = 0;rain_draw[62][125] = 0;rain_draw[63][125] = 0;rain_draw[64][125] = 0;rain_draw[65][125] = 0;rain_draw[66][125] = 0;rain_draw[67][125] = 0;rain_draw[68][125] = 0;rain_draw[69][125] = 0;rain_draw[70][125] = 0;rain_draw[71][125] = 0;rain_draw[72][125] = 0;rain_draw[73][125] = 0;rain_draw[74][125] = 0;rain_draw[75][125] = 0;rain_draw[76][125] = 0;rain_draw[77][125] = 0;rain_draw[78][125] = 0;rain_draw[79][125] = 0;rain_draw[80][125] = 0;rain_draw[81][125] = 0;rain_draw[82][125] = 0;rain_draw[83][125] = 0;rain_draw[84][125] = 0;rain_draw[85][125] = 0;rain_draw[86][125] = 0;rain_draw[87][125] = 0;rain_draw[88][125] = 0;rain_draw[89][125] = 0;rain_draw[90][125] = 0;rain_draw[91][125] = 0;rain_draw[92][125] = 0;rain_draw[93][125] = 0;rain_draw[94][125] = 0;rain_draw[95][125] = 0;
        rain_draw[0][126] = 0;rain_draw[1][126] = 0;rain_draw[2][126] = 0;rain_draw[3][126] = 0;rain_draw[4][126] = 0;rain_draw[5][126] = 0;rain_draw[6][126] = 0;rain_draw[7][126] = 0;rain_draw[8][126] = 0;rain_draw[9][126] = 0;rain_draw[10][126] = 0;rain_draw[11][126] = 0;rain_draw[12][126] = 0;rain_draw[13][126] = 0;rain_draw[14][126] = 0;rain_draw[15][126] = 0;rain_draw[16][126] = 0;rain_draw[17][126] = 0;rain_draw[18][126] = 0;rain_draw[19][126] = 0;rain_draw[20][126] = 0;rain_draw[21][126] = 0;rain_draw[22][126] = 0;rain_draw[23][126] = 0;rain_draw[24][126] = 0;rain_draw[25][126] = 0;rain_draw[26][126] = 0;rain_draw[27][126] = 0;rain_draw[28][126] = 0;rain_draw[29][126] = 0;rain_draw[30][126] = 0;rain_draw[31][126] = 0;rain_draw[32][126] = 0;rain_draw[33][126] = 0;rain_draw[34][126] = 0;rain_draw[35][126] = 0;rain_draw[36][126] = 0;rain_draw[37][126] = 0;rain_draw[38][126] = 0;rain_draw[39][126] = 0;rain_draw[40][126] = 0;rain_draw[41][126] = 0;rain_draw[42][126] = 0;rain_draw[43][126] = 0;rain_draw[44][126] = 0;rain_draw[45][126] = 0;rain_draw[46][126] = 0;rain_draw[47][126] = 0;rain_draw[48][126] = 0;rain_draw[49][126] = 0;rain_draw[50][126] = 0;rain_draw[51][126] = 0;rain_draw[52][126] = 0;rain_draw[53][126] = 0;rain_draw[54][126] = 0;rain_draw[55][126] = 0;rain_draw[56][126] = 0;rain_draw[57][126] = 0;rain_draw[58][126] = 0;rain_draw[59][126] = 0;rain_draw[60][126] = 0;rain_draw[61][126] = 0;rain_draw[62][126] = 0;rain_draw[63][126] = 0;rain_draw[64][126] = 0;rain_draw[65][126] = 0;rain_draw[66][126] = 0;rain_draw[67][126] = 0;rain_draw[68][126] = 0;rain_draw[69][126] = 0;rain_draw[70][126] = 0;rain_draw[71][126] = 0;rain_draw[72][126] = 0;rain_draw[73][126] = 0;rain_draw[74][126] = 0;rain_draw[75][126] = 0;rain_draw[76][126] = 0;rain_draw[77][126] = 0;rain_draw[78][126] = 0;rain_draw[79][126] = 0;rain_draw[80][126] = 0;rain_draw[81][126] = 0;rain_draw[82][126] = 0;rain_draw[83][126] = 0;rain_draw[84][126] = 0;rain_draw[85][126] = 0;rain_draw[86][126] = 0;rain_draw[87][126] = 0;rain_draw[88][126] = 0;rain_draw[89][126] = 0;rain_draw[90][126] = 0;rain_draw[91][126] = 0;rain_draw[92][126] = 0;rain_draw[93][126] = 0;rain_draw[94][126] = 0;rain_draw[95][126] = 0;
        rain_draw[0][127] = 0;rain_draw[1][127] = 0;rain_draw[2][127] = 0;rain_draw[3][127] = 0;rain_draw[4][127] = 0;rain_draw[5][127] = 0;rain_draw[6][127] = 0;rain_draw[7][127] = 0;rain_draw[8][127] = 0;rain_draw[9][127] = 0;rain_draw[10][127] = 0;rain_draw[11][127] = 0;rain_draw[12][127] = 0;rain_draw[13][127] = 0;rain_draw[14][127] = 0;rain_draw[15][127] = 0;rain_draw[16][127] = 0;rain_draw[17][127] = 0;rain_draw[18][127] = 0;rain_draw[19][127] = 0;rain_draw[20][127] = 0;rain_draw[21][127] = 0;rain_draw[22][127] = 0;rain_draw[23][127] = 0;rain_draw[24][127] = 0;rain_draw[25][127] = 0;rain_draw[26][127] = 0;rain_draw[27][127] = 0;rain_draw[28][127] = 0;rain_draw[29][127] = 0;rain_draw[30][127] = 0;rain_draw[31][127] = 0;rain_draw[32][127] = 0;rain_draw[33][127] = 0;rain_draw[34][127] = 0;rain_draw[35][127] = 0;rain_draw[36][127] = 0;rain_draw[37][127] = 0;rain_draw[38][127] = 0;rain_draw[39][127] = 0;rain_draw[40][127] = 0;rain_draw[41][127] = 0;rain_draw[42][127] = 0;rain_draw[43][127] = 0;rain_draw[44][127] = 0;rain_draw[45][127] = 0;rain_draw[46][127] = 0;rain_draw[47][127] = 0;rain_draw[48][127] = 0;rain_draw[49][127] = 0;rain_draw[50][127] = 0;rain_draw[51][127] = 0;rain_draw[52][127] = 0;rain_draw[53][127] = 0;rain_draw[54][127] = 0;rain_draw[55][127] = 0;rain_draw[56][127] = 0;rain_draw[57][127] = 0;rain_draw[58][127] = 0;rain_draw[59][127] = 0;rain_draw[60][127] = 0;rain_draw[61][127] = 0;rain_draw[62][127] = 0;rain_draw[63][127] = 0;rain_draw[64][127] = 0;rain_draw[65][127] = 0;rain_draw[66][127] = 0;rain_draw[67][127] = 0;rain_draw[68][127] = 0;rain_draw[69][127] = 0;rain_draw[70][127] = 0;rain_draw[71][127] = 0;rain_draw[72][127] = 0;rain_draw[73][127] = 0;rain_draw[74][127] = 0;rain_draw[75][127] = 0;rain_draw[76][127] = 0;rain_draw[77][127] = 0;rain_draw[78][127] = 0;rain_draw[79][127] = 0;rain_draw[80][127] = 0;rain_draw[81][127] = 0;rain_draw[82][127] = 0;rain_draw[83][127] = 0;rain_draw[84][127] = 0;rain_draw[85][127] = 0;rain_draw[86][127] = 0;rain_draw[87][127] = 0;rain_draw[88][127] = 0;rain_draw[89][127] = 0;rain_draw[90][127] = 0;rain_draw[91][127] = 0;rain_draw[92][127] = 0;rain_draw[93][127] = 0;rain_draw[94][127] = 0;rain_draw[95][127] = 0;
    end

    
end


assign active_rain = (rain_draw[v_counter][h_counter]) ? 1 : 0;


endmodule